`timescale 1ns / 1ps
module gameO_214x160_rom(
    input  [7:0] x_idx,
    input  [7:0] y_idx,
    output reg [7:0] RED,
    output reg [7:0] GRN,
    output reg [7:0] BLU);
always @ (*)
    case ({y_idx,x_idx})
        0:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        41:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        42:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        43:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        44:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        45:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        46:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        47:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        48:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        49:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        50:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        51:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        52:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        53:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        54:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        55:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        56:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        57:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        58:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        59:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        60:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        61:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        62:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        63:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        64:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        65:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        66:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        67:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        68:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        69:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        70:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        71:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        72:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        73:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        74:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        75:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        76:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        77:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        78:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        79:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        80:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        81:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        82:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        83:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        84:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        85:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        86:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        87:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        88:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        89:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        90:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        91:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        92:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        93:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        94:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        95:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        96:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        97:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        98:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        99:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8463:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd16;
        end
        8464:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd25;
        end
        8465:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd22;
        end
        8466:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        8467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8574:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd17;
        end
        8575:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd25;
        end
        8576:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd25;
        end
        8577:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd17;
        end
        8578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8716:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd4;
        end
        8717:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd62;
        end
        8718:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd92;
        end
        8719:
        begin
            RED=8'd0;
            GRN=8'd79;
            BLU=8'd114;
        end
        8720:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd125;
        end
        8721:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd121;
        end
        8722:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd94;
        end
        8723:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd68;
        end
        8724:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd8;
        end
        8725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8740:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd18;
        end
        8741:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8742:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8743:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8744:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8745:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8746:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8747:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd13;
        end
        8748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8756:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd5;
        end
        8757:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8758:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8759:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8760:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8761:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8762:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8763:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8764:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8765:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd2;
        end
        8766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8773:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd13;
        end
        8774:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8775:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8776:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8777:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8778:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8779:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8780:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8781:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8782:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd2;
        end
        8783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd6;
        end
        8787:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd21;
        end
        8788:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8789:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8790:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8791:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8792:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8793:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8794:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8795:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8796:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8797:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8798:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8799:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8800:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8801:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8802:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8803:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8804:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd12;
        end
        8805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8827:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd6;
        end
        8828:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd65;
        end
        8829:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd93;
        end
        8830:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd115;
        end
        8831:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd125;
        end
        8832:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd125;
        end
        8833:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd114;
        end
        8834:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd87;
        end
        8835:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd53;
        end
        8836:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd3;
        end
        8837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8844:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd12;
        end
        8845:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8846:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8847:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8848:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8849:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8850:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8851:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8852:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd16;
        end
        8853:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        8854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8863:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd18;
        end
        8864:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8865:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8866:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd19;
        end
        8867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd9;
        end
        8869:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8870:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8871:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8872:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8873:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8874:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8875:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8876:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8877:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8878:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8879:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8880:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8881:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8882:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8883:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8884:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8885:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8886:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd9;
        end
        8887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8890:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd18;
        end
        8891:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8892:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8893:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8894:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8895:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8896:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8897:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8898:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8899:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8900:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8901:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8902:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd21;
        end
        8903:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd10;
        end
        8904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8971:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd15;
        end
        8972:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd77;
        end
        8973:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd179;
        end
        8974:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd229;
        end
        8975:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        8976:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        8977:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        8978:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        8979:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd188;
        end
        8980:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd83;
        end
        8981:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd18;
        end
        8982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8995:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd11;
        end
        8996:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd100;
        end
        8997:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        8998:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        8999:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9000:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9001:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9002:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9003:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd76;
        end
        9004:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        9005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9012:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd32;
        end
        9013:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd110;
        end
        9014:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9015:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9016:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9017:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9018:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9019:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9020:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9021:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd31;
        end
        9022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9029:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd67;
        end
        9030:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9031:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9032:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9033:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9034:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9035:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9036:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9037:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9038:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd13;
        end
        9039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9042:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd31;
        end
        9043:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd109;
        end
        9044:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9045:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9046:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9047:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9048:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9049:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9050:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9051:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9052:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9053:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9054:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9055:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9056:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9057:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9058:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9059:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9060:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd68;
        end
        9061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9082:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd25;
        end
        9083:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd86;
        end
        9084:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd183;
        end
        9085:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd230;
        end
        9086:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9087:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9088:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9089:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9090:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd220;
        end
        9091:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd163;
        end
        9092:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd74;
        end
        9093:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd12;
        end
        9094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9100:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd52;
        end
        9101:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9102:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9103:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9104:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9105:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9106:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9107:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9108:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd100;
        end
        9109:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd11;
        end
        9110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd8;
        end
        9119:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd98;
        end
        9120:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9121:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9122:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd89;
        end
        9123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9124:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd45;
        end
        9125:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9126:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9127:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9128:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9129:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9130:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9131:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9132:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9133:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9134:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9135:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9136:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9137:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9138:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9139:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9140:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9141:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9142:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd53;
        end
        9143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9146:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd89;
        end
        9147:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9148:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9149:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9150:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9151:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9152:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9153:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9154:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9155:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9156:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9157:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9158:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd110;
        end
        9159:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd91;
        end
        9160:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd72;
        end
        9161:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd43;
        end
        9162:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd6;
        end
        9163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9226:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd13;
        end
        9227:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd89;
        end
        9228:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd218;
        end
        9229:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9230:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9231:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9232:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9233:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9234:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9235:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9236:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd220;
        end
        9237:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd91;
        end
        9238:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd6;
        end
        9239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9251:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd36;
        end
        9252:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd218;
        end
        9253:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9254:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9255:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9256:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9257:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9258:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9259:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd170;
        end
        9260:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd2;
        end
        9261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9268:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        9269:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        9270:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9271:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9272:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9273:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9274:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9275:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9276:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9277:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd95;
        end
        9278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9285:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd150;
        end
        9286:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9287:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9288:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9289:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9290:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9291:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9292:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9293:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9294:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        9295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9298:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        9299:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        9300:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9301:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9302:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9303:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9304:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9305:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9306:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9307:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9308:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9309:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9310:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9311:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9312:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9313:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9314:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9315:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9316:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd151;
        end
        9317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9337:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd21;
        end
        9338:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd113;
        end
        9339:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd232;
        end
        9340:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9341:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9342:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9343:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9344:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9345:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9347:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9348:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd219;
        end
        9349:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd80;
        end
        9350:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd9;
        end
        9351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9356:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd96;
        end
        9357:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9358:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9359:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9360:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9361:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9362:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9363:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9364:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd226;
        end
        9365:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd42;
        end
        9366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9374:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd27;
        end
        9375:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd212;
        end
        9376:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9377:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9378:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd171;
        end
        9379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9380:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        9381:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9382:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9383:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9384:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9385:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9386:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9387:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9388:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9389:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9390:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9391:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9393:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9394:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9396:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9397:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9398:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd119;
        end
        9399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9402:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        9403:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9404:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9405:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9406:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9407:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9408:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9409:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9410:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9411:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9412:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9413:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9414:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9415:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9416:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd224;
        end
        9417:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd158;
        end
        9418:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd67;
        end
        9419:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd13;
        end
        9420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        9482:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd78;
        end
        9483:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd220;
        end
        9484:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9485:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9486:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9487:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9488:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9489:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9490:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9491:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9492:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9493:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd210;
        end
        9494:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd46;
        end
        9495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9507:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd47;
        end
        9508:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd224;
        end
        9509:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9510:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9511:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9512:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9513:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9514:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9515:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd185;
        end
        9516:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd5;
        end
        9517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9524:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        9525:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        9526:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9527:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9528:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9529:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9530:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9531:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9532:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9533:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd122;
        end
        9534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        9541:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd182;
        end
        9542:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9543:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9544:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9545:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9546:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9547:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9548:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9549:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9550:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        9551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9554:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        9555:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        9556:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9557:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9558:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9559:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9560:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9561:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9562:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9563:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9564:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9565:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9566:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9567:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9568:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9569:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9570:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9571:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9572:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd151;
        end
        9573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9592:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd9;
        end
        9593:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd109;
        end
        9594:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd228;
        end
        9595:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9596:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9597:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9598:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9599:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9600:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9601:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9603:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9604:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9605:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd221;
        end
        9606:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd62;
        end
        9607:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd1;
        end
        9608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9612:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd80;
        end
        9613:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        9614:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9615:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9616:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9617:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9618:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9619:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9620:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9621:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd68;
        end
        9622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9630:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd38;
        end
        9631:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd219;
        end
        9632:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9633:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9634:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd143;
        end
        9635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9636:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        9637:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9638:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9639:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9640:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9641:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9642:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9643:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9644:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9645:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9646:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9647:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9648:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9649:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9650:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9652:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9653:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9654:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd119;
        end
        9655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9658:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        9659:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9660:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9661:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9662:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9663:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9664:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9665:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9666:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9667:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9668:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9669:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9670:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9671:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9673:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9674:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd220;
        end
        9675:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd83;
        end
        9676:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd10;
        end
        9677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9737:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd16;
        end
        9738:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd208;
        end
        9739:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9740:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9741:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9742:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9743:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9744:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9745:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9746:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9747:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9748:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9749:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9750:
        begin
            RED=8'd0;
            GRN=8'd122;
            BLU=8'd161;
        end
        9751:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd4;
        end
        9752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9763:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd64;
        end
        9764:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd232;
        end
        9765:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9766:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9767:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9768:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9769:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9770:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9771:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd210;
        end
        9772:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd8;
        end
        9773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9780:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        9781:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        9782:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9783:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9784:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9785:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9786:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9787:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9788:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9789:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd155;
        end
        9790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9796:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd4;
        end
        9797:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd208;
        end
        9798:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9799:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9800:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9801:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9802:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9803:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9804:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9805:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9806:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        9807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9810:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        9811:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        9812:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9813:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9814:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9815:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9816:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9817:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9818:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9819:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9820:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9821:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9822:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9823:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9824:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9825:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9826:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9827:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9828:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd151;
        end
        9829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9848:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd65;
        end
        9849:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd222;
        end
        9850:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9851:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9852:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9853:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9854:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9855:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9856:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9857:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9859:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9860:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9861:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9862:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd198;
        end
        9863:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd15;
        end
        9864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9868:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd51;
        end
        9869:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd231;
        end
        9870:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9871:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9872:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9873:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9874:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9875:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9876:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9877:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd96;
        end
        9878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9886:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd55;
        end
        9887:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd227;
        end
        9888:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9889:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9890:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd109;
        end
        9891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9892:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        9893:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9894:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9895:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9896:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9897:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9898:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9899:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9900:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9901:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9902:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9903:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9904:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9905:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9906:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9908:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9909:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9910:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd119;
        end
        9911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9914:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        9915:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9916:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9917:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9918:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9919:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9920:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9921:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9922:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9923:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9924:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9925:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9926:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9927:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9928:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9929:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9930:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9932:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd72;
        end
        9933:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd2;
        end
        9934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9993:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd141;
        end
        9994:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9995:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9996:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9997:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9998:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        9999:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10000:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10001:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10002:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10003:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10004:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10005:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10006:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd222;
        end
        10007:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd45;
        end
        10008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10019:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd100;
        end
        10020:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10021:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10022:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10023:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10024:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10025:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10026:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10027:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10028:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd11;
        end
        10029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10036:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        10037:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        10038:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10039:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10040:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10041:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10042:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10043:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10044:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10045:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd170;
        end
        10046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10052:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd5;
        end
        10053:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd232;
        end
        10054:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10055:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10056:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10057:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10058:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10059:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10060:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10061:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10062:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        10063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10066:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        10067:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        10068:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10069:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10070:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10071:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10072:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10073:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10074:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10075:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10076:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10077:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10078:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10079:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10080:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10081:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10082:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10083:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10084:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd151;
        end
        10085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10104:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd184;
        end
        10105:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10106:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10107:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10108:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10109:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10110:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10113:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10114:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10115:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10116:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10117:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10118:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10119:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd116;
        end
        10120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10124:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd27;
        end
        10125:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd223;
        end
        10126:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10127:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10128:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10129:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10130:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10131:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10132:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10133:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd110;
        end
        10134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10142:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd83;
        end
        10143:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd232;
        end
        10144:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10145:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10146:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd97;
        end
        10147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10148:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        10149:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10150:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10151:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10152:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10153:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10154:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10155:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10156:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10157:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10158:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10159:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10161:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10162:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10164:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10165:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10166:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd119;
        end
        10167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10170:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        10171:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10172:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10173:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10174:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10175:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10176:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10177:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10178:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10179:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10180:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10181:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10182:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10183:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10185:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10186:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10188:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd212;
        end
        10189:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd25;
        end
        10190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10248:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd45;
        end
        10249:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd223;
        end
        10250:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10251:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10252:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10253:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10254:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10255:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10256:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10257:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10258:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10259:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10260:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10261:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10262:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10263:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd132;
        end
        10264:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd0;
        end
        10265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10275:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd130;
        end
        10276:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10277:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10278:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10279:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10280:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10281:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10282:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10283:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10284:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd32;
        end
        10285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10292:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        10293:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        10294:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10295:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10296:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10297:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10298:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10299:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10300:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10301:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd199;
        end
        10302:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd0;
        end
        10303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10308:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd27;
        end
        10309:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd232;
        end
        10310:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10311:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10312:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10313:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10314:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10315:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10316:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10317:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10318:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        10319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10322:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        10323:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        10324:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10325:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10326:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10327:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10328:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10329:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10330:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10331:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10332:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10333:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10334:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10335:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10336:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10337:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10338:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10339:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10340:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd151;
        end
        10341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10359:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd97;
        end
        10360:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        10361:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10362:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10363:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10364:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10365:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10366:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd215;
        end
        10367:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd48;
        end
        10368:
        begin
            RED=8'd0;
            GRN=8'd82;
            BLU=8'd133;
        end
        10369:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10370:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10371:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10372:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10373:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10374:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10375:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd215;
        end
        10376:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd27;
        end
        10377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10380:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd22;
        end
        10381:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd213;
        end
        10382:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10383:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10384:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10385:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10386:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10387:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10388:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10389:
        begin
            RED=8'd0;
            GRN=8'd122;
            BLU=8'd137;
        end
        10390:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        10391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10398:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd116;
        end
        10399:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10400:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10401:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10402:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd68;
        end
        10403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10404:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        10405:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10406:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10407:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10408:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10409:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10410:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10411:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10412:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10413:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10414:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10415:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10417:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10418:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10420:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10421:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10422:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd119;
        end
        10423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10426:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        10427:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10428:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10429:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10430:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10431:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10432:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10433:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10434:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10435:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10436:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10437:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10438:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10439:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10441:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10442:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10443:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10444:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10445:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd147;
        end
        10446:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd0;
        end
        10447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10504:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd139;
        end
        10505:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd231;
        end
        10506:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10507:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10508:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10509:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10510:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10511:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10512:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd130;
        end
        10513:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd27;
        end
        10514:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd113;
        end
        10515:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd225;
        end
        10516:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10517:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10518:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10519:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd204;
        end
        10520:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd16;
        end
        10521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10531:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd156;
        end
        10532:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10533:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10534:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10535:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10536:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10537:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10538:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10539:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10540:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd62;
        end
        10541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10548:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        10549:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        10550:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10551:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10552:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10553:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10554:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10555:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10556:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10557:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd215;
        end
        10558:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd16;
        end
        10559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10564:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd56;
        end
        10565:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        10566:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10567:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10568:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10569:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10570:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10571:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10572:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10573:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10574:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        10575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10578:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        10579:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        10580:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10581:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10582:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10583:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10584:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10585:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10586:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10587:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10588:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10589:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10590:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10591:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10592:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10593:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10594:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10595:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10596:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd151;
        end
        10597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd14;
        end
        10615:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd188;
        end
        10616:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10617:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10618:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10619:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10620:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10621:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10622:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd105;
        end
        10623:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd4;
        end
        10624:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd20;
        end
        10625:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd193;
        end
        10626:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10627:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10628:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10629:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10630:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10631:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd230;
        end
        10632:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd114;
        end
        10633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10636:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd13;
        end
        10637:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd195;
        end
        10638:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10639:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10640:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10641:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10642:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10643:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10644:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10645:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd157;
        end
        10646:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        10647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10654:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd130;
        end
        10655:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10656:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10657:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10658:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd38;
        end
        10659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10660:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        10661:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10662:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10663:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10664:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10665:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10666:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10667:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10668:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10669:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10670:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10671:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10673:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10674:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10676:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10677:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10678:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd119;
        end
        10679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10682:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        10683:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10684:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10685:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10686:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10687:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10688:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10689:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10690:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10691:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10692:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10693:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10694:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10695:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10696:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10698:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10699:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10700:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10701:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd225;
        end
        10702:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd42;
        end
        10703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10759:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd39;
        end
        10760:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd218;
        end
        10761:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10762:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10763:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10764:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10765:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10766:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10767:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd156;
        end
        10768:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd20;
        end
        10769:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd1;
        end
        10770:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd17;
        end
        10771:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd105;
        end
        10772:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10773:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10774:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10775:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        10776:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd67;
        end
        10777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        10787:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd171;
        end
        10788:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10789:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10790:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10791:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10792:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10793:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10794:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10795:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10796:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd89;
        end
        10797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10804:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        10805:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        10806:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10807:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10808:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10809:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10810:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10811:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10812:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10813:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd219;
        end
        10814:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd29;
        end
        10815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10820:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd83;
        end
        10821:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10822:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10823:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10824:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10825:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10826:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10827:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10828:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10829:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10830:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        10831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10834:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        10835:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        10836:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10837:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10838:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10839:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10840:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10841:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10842:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10843:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd83;
        end
        10844:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10845:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10846:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10847:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10848:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10849:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10850:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10851:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10852:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd24;
        end
        10853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10870:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd65;
        end
        10871:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd226;
        end
        10872:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10873:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10874:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10875:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10876:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10877:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd218;
        end
        10878:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd30;
        end
        10879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        10881:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd118;
        end
        10882:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        10883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10884:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10885:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10886:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10887:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10888:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd181;
        end
        10889:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd10;
        end
        10890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd8;
        end
        10893:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd183;
        end
        10894:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10895:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10896:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10897:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10898:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10899:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10900:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10901:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd185;
        end
        10902:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        10903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10910:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd153;
        end
        10911:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10912:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10913:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd223;
        end
        10914:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd16;
        end
        10915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10916:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        10917:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10918:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10919:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10920:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10921:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10922:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10923:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10924:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd220;
        end
        10925:
        begin
            RED=8'd0;
            GRN=8'd59;
            BLU=8'd68;
        end
        10926:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10927:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10928:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10929:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10930:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10931:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10932:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10933:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10934:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd19;
        end
        10935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10938:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        10939:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10940:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10941:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10942:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10943:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10944:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10945:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10946:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd174;
        end
        10947:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd38;
        end
        10948:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd78;
        end
        10949:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd199;
        end
        10950:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10951:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10952:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10954:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10955:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10956:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10957:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        10958:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd126;
        end
        10959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11015:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd103;
        end
        11016:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        11017:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11018:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11019:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11020:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11021:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11022:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd227;
        end
        11023:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd49;
        end
        11024:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        11025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11027:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd24;
        end
        11028:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd194;
        end
        11029:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11030:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11031:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11032:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd125;
        end
        11033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11042:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd10;
        end
        11043:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd193;
        end
        11044:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11045:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11046:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11047:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11048:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11049:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11050:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11051:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11052:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd104;
        end
        11053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11060:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        11061:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        11062:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11063:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11064:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11065:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11066:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11067:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11068:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11069:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd224;
        end
        11070:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd49;
        end
        11071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11076:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd98;
        end
        11077:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11078:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11079:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11080:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11081:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11082:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11083:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11084:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11085:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11086:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        11087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11090:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        11091:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        11092:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11093:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11094:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11095:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11096:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11097:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11098:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11099:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        11100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11126:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd135;
        end
        11127:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        11128:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11129:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11130:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11131:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11132:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11133:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd179;
        end
        11134:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd4;
        end
        11135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11137:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd60;
        end
        11138:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd227;
        end
        11139:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11140:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11141:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11142:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11143:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11144:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd222;
        end
        11145:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd41;
        end
        11146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        11149:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd160;
        end
        11150:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11151:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11152:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11153:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11154:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11155:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11156:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11157:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd201;
        end
        11158:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        11159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd7;
        end
        11166:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd181;
        end
        11167:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11168:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11169:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd211;
        end
        11170:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd10;
        end
        11171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11172:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        11173:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11174:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11175:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11176:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11177:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11178:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11179:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11180:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        11181:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        11182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11194:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        11195:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11196:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11197:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11198:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11199:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11200:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11201:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11202:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        11203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11204:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd12;
        end
        11205:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd61;
        end
        11206:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd210;
        end
        11207:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11208:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11210:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11211:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11212:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11213:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11214:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd199;
        end
        11215:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd0;
        end
        11216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11271:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd177;
        end
        11272:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11273:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11274:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11275:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11276:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11277:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11278:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd173;
        end
        11279:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd6;
        end
        11280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11283:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd2;
        end
        11284:
        begin
            RED=8'd0;
            GRN=8'd73;
            BLU=8'd131;
        end
        11285:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11286:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11287:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11288:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd173;
        end
        11289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11298:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd17;
        end
        11299:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd215;
        end
        11300:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11301:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11302:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11303:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11304:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11305:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11306:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11307:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11308:
        begin
            RED=8'd0;
            GRN=8'd116;
            BLU=8'd133;
        end
        11309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11316:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        11317:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        11318:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11319:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11320:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11321:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11322:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11323:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11324:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11325:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        11326:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd70;
        end
        11327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11332:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd127;
        end
        11333:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11334:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11335:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11336:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11337:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11338:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11339:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11340:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11341:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11342:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        11343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11346:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        11347:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        11348:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11349:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11350:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11351:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11352:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11353:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11354:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11355:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        11356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11382:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd196;
        end
        11383:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11384:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11385:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11386:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11387:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11388:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11389:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd131;
        end
        11390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11393:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd15;
        end
        11394:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd221;
        end
        11395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11396:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11397:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11398:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11399:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11400:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11401:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd102;
        end
        11402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11405:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd133;
        end
        11406:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11407:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11408:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11409:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11410:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11411:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11412:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11413:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd223;
        end
        11414:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd2;
        end
        11415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11421:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd14;
        end
        11422:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd203;
        end
        11423:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11424:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11425:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd190;
        end
        11426:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd6;
        end
        11427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11428:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        11429:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11430:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11431:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11432:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11433:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11434:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11435:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11436:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        11437:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        11438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11450:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        11451:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11452:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11453:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11454:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11455:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11456:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11457:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11458:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        11459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11461:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd6;
        end
        11462:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd139;
        end
        11463:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        11464:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11465:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11466:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11467:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11468:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11469:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11470:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        11471:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd39;
        end
        11472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11526:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd34;
        end
        11527:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd218;
        end
        11528:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11529:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11530:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11531:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11532:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11533:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11534:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd110;
        end
        11535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11540:
        begin
            RED=8'd0;
            GRN=8'd33;
            BLU=8'd70;
        end
        11541:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd228;
        end
        11542:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11543:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11544:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd207;
        end
        11545:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd11;
        end
        11546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11554:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd34;
        end
        11555:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd228;
        end
        11556:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11557:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11558:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11559:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11560:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11561:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11562:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11563:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11564:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd164;
        end
        11565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11572:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        11573:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        11574:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11575:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11576:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11577:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11578:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11579:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11580:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11581:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11582:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd99;
        end
        11583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11588:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd158;
        end
        11589:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11590:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11591:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11592:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11593:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11594:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11595:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11596:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11597:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11598:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        11599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11602:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        11603:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        11604:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11605:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11606:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11607:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11608:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11609:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11610:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11611:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        11612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11637:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd40;
        end
        11638:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd225;
        end
        11639:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11640:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11641:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11642:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11643:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11644:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11645:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd89;
        end
        11646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11650:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd192;
        end
        11651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11652:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11653:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11654:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11655:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11656:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11657:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd167;
        end
        11658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11661:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd115;
        end
        11662:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11663:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11664:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11665:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11666:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11667:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11668:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11669:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11670:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd25;
        end
        11671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11677:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd18;
        end
        11678:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd218;
        end
        11679:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11680:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11681:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd162;
        end
        11682:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd2;
        end
        11683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11684:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        11685:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11686:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11687:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11688:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11689:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11690:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11691:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11692:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        11693:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        11694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11706:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        11707:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11708:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11709:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11710:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11711:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11712:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11713:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11714:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        11715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11718:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd55;
        end
        11719:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd228;
        end
        11720:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11721:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11722:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11723:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11724:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11725:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11726:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        11727:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd95;
        end
        11728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11782:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd98;
        end
        11783:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd230;
        end
        11784:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11785:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11786:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11787:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11788:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11789:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11790:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd56;
        end
        11791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11796:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd33;
        end
        11797:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd215;
        end
        11798:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11799:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11800:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd224;
        end
        11801:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd39;
        end
        11802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11810:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd60;
        end
        11811:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        11812:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11813:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11814:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11815:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11816:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11817:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11818:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11819:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11820:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd183;
        end
        11821:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd0;
        end
        11822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11828:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        11829:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        11830:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11831:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11832:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11833:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11834:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11835:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11836:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11837:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11838:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd123;
        end
        11839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11844:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd184;
        end
        11845:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11846:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11847:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11848:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11849:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11850:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11851:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11852:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11853:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11854:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        11855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11858:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        11859:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        11860:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11861:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11862:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11863:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11864:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11865:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11866:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11867:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        11868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11893:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd92;
        end
        11894:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd231;
        end
        11895:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11896:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11897:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11898:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11899:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11900:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11901:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd64;
        end
        11902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11906:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd158;
        end
        11907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11908:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11909:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11910:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11911:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11912:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11913:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd210;
        end
        11914:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd10;
        end
        11915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11917:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd89;
        end
        11918:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd232;
        end
        11919:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11920:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11921:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11922:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11923:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11924:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11925:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11926:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd48;
        end
        11927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11933:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd32;
        end
        11934:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd227;
        end
        11935:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11936:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11937:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd135;
        end
        11938:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        11939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11940:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        11941:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11942:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11943:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11944:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11945:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11946:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11947:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11948:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        11949:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        11950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11962:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        11963:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11964:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11965:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11966:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11967:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11968:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11969:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11970:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        11971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd9;
        end
        11975:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd202;
        end
        11976:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11977:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11978:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11979:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11980:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11981:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11982:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        11983:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd136;
        end
        11984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        12038:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd159;
        end
        12039:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12040:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12041:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12042:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12043:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12044:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12045:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd219;
        end
        12046:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd24;
        end
        12047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd12;
        end
        12053:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd197;
        end
        12054:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12055:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12056:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        12057:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd77;
        end
        12058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12066:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd82;
        end
        12067:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12068:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12069:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12070:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12071:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12072:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12073:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12074:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12075:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12076:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd199;
        end
        12077:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd6;
        end
        12078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12084:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        12085:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        12086:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12087:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12088:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12089:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12090:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12091:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12092:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12093:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12094:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd143;
        end
        12095:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        12096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd6;
        end
        12100:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd201;
        end
        12101:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12102:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12103:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12104:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12105:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12106:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12107:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12108:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12109:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12110:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        12111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12114:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        12115:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        12116:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12117:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12118:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12119:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12120:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12121:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12122:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12123:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        12124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12149:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd142;
        end
        12150:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12151:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12152:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12153:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12154:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12155:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12156:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12157:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd40;
        end
        12158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12162:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd133;
        end
        12163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12164:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12165:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12166:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12167:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12168:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12169:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd227;
        end
        12170:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd43;
        end
        12171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12173:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd66;
        end
        12174:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd230;
        end
        12175:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12176:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12177:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12178:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12179:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12180:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12181:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12182:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd69;
        end
        12183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12189:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd58;
        end
        12190:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        12191:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12192:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12193:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd115;
        end
        12194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12196:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        12197:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12198:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12199:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12200:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12201:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12202:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12203:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12204:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        12205:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        12206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12218:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        12219:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12220:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12221:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12222:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12223:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12224:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12225:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12226:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        12227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12231:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd166;
        end
        12232:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12233:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12234:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12235:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12236:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12237:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12238:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12239:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd168;
        end
        12240:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd4;
        end
        12241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12293:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd19;
        end
        12294:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd202;
        end
        12295:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12296:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12297:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12298:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12299:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12300:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12301:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd195;
        end
        12302:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd13;
        end
        12303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12309:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd178;
        end
        12310:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12311:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12312:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12313:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd113;
        end
        12314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12322:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd100;
        end
        12323:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12324:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12325:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12326:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12327:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12328:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12329:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12330:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12331:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12332:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd213;
        end
        12333:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd23;
        end
        12334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12340:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        12341:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        12342:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12343:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12344:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12345:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12347:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12348:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12349:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12350:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd169;
        end
        12351:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd3;
        end
        12352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12355:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd21;
        end
        12356:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd209;
        end
        12357:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12358:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12359:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12360:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12361:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12362:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12363:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12364:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12365:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12366:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        12367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12370:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        12371:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        12372:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12373:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12374:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12375:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12376:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12377:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12378:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12379:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        12380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd8;
        end
        12405:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd188;
        end
        12406:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12407:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12408:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12409:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12410:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12411:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12412:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        12413:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd17;
        end
        12414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12418:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd116;
        end
        12419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12420:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12421:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12422:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12423:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12424:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12425:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        12426:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd92;
        end
        12427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12429:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd53;
        end
        12430:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd225;
        end
        12431:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12432:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12433:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12434:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12435:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12436:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12437:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12438:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd89;
        end
        12439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12445:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd82;
        end
        12446:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12447:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12448:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12449:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd95;
        end
        12450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12452:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        12453:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12454:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12455:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12456:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12457:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12458:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12459:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12460:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        12461:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        12462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12474:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        12475:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12476:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12477:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12478:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12479:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12480:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12481:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12482:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        12483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12487:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd135;
        end
        12488:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12489:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12490:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12491:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12492:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12493:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12494:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12495:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd193;
        end
        12496:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd12;
        end
        12497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12549:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd49;
        end
        12550:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd227;
        end
        12551:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12552:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12553:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12554:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12555:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12556:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12557:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd176;
        end
        12558:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd5;
        end
        12559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12565:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd156;
        end
        12566:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12567:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12568:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12569:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd143;
        end
        12570:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        12571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12578:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd128;
        end
        12579:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12580:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12581:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12582:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12583:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12584:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12585:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12586:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12587:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12588:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd221;
        end
        12589:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd41;
        end
        12590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12596:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        12597:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        12598:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12599:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12600:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12601:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12603:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12604:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12605:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12606:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd191;
        end
        12607:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd11;
        end
        12608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12611:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd40;
        end
        12612:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd220;
        end
        12613:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12614:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12615:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12616:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12617:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12618:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12619:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12620:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12621:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12622:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        12623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12626:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        12627:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        12628:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12629:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12630:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12631:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12632:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12633:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12634:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12635:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        12636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12660:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd27;
        end
        12661:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd211;
        end
        12662:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12663:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12664:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12665:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12666:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12667:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12668:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd218;
        end
        12669:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd14;
        end
        12670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12674:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd104;
        end
        12675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12676:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12677:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12678:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12679:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12680:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12681:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12682:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd133;
        end
        12683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12685:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd33;
        end
        12686:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd218;
        end
        12687:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12688:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12689:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12690:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12691:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12692:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12693:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12694:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd108;
        end
        12695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12701:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd99;
        end
        12702:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12703:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12704:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        12705:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd66;
        end
        12706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12708:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        12709:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12710:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12711:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12712:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12713:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12714:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12715:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12716:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        12717:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        12718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12730:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        12731:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12732:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12733:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12734:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12735:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12736:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12737:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12738:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        12739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12743:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd105;
        end
        12744:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12745:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12746:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12747:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12748:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12749:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12750:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12751:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd202;
        end
        12752:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd19;
        end
        12753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12805:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd89;
        end
        12806:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12807:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12808:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12809:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12810:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12811:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12812:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12813:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd160;
        end
        12814:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd0;
        end
        12815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12821:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd142;
        end
        12822:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12823:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12824:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12825:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd169;
        end
        12826:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd2;
        end
        12827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12834:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd163;
        end
        12835:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12836:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12837:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12838:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12839:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12840:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12841:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12842:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12843:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12844:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd225;
        end
        12845:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd52;
        end
        12846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12852:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        12853:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        12854:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12855:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12856:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12857:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12859:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12860:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12861:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12862:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd208;
        end
        12863:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd22;
        end
        12864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12867:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd55;
        end
        12868:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd228;
        end
        12869:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12870:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12871:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12872:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12873:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12874:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12875:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12876:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12877:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12878:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        12879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12882:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        12883:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        12884:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12885:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12886:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12887:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12888:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12889:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12890:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12891:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        12892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12916:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd46;
        end
        12917:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd222;
        end
        12918:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12919:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12920:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12921:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12922:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12923:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12924:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd207;
        end
        12925:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd12;
        end
        12926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12930:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd91;
        end
        12931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12932:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12933:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12934:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12935:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12936:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12937:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12938:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd162;
        end
        12939:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd2;
        end
        12940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd13;
        end
        12942:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd211;
        end
        12943:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12944:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12945:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12946:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12947:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12948:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12949:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12950:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd140;
        end
        12951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12957:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd126;
        end
        12958:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12959:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12960:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd223;
        end
        12961:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd42;
        end
        12962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12964:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        12965:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12966:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12967:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12968:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12969:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12970:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12971:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12972:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        12973:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        12974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12986:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        12987:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12988:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12989:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12990:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12991:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12992:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12993:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        12994:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        12995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        12999:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd84;
        end
        13000:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13001:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13002:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13003:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13004:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13005:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13006:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13007:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd210;
        end
        13008:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd25;
        end
        13009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13061:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd130;
        end
        13062:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13063:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13064:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13065:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13066:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13067:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13068:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13069:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd136;
        end
        13070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13077:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd130;
        end
        13078:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13079:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13080:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13081:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd190;
        end
        13082:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd10;
        end
        13083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13090:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd189;
        end
        13091:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13092:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13093:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13094:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13095:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13096:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13097:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13098:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13099:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13100:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13101:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd72;
        end
        13102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13108:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        13109:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        13110:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13113:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13114:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13115:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13116:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13117:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13118:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd217;
        end
        13119:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd28;
        end
        13120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13123:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd66;
        end
        13124:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd232;
        end
        13125:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13126:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13127:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13128:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13129:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13130:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13131:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13132:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13133:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13134:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        13135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13138:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        13139:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        13140:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13141:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13142:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13143:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13144:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13145:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13146:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13147:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        13148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13172:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd80;
        end
        13173:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        13174:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13175:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13176:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13177:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13178:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13179:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13180:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd195;
        end
        13181:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd10;
        end
        13182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13186:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd77;
        end
        13187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13188:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13189:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13190:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13191:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13192:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13193:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13194:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd196;
        end
        13195:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd13;
        end
        13196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13198:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd203;
        end
        13199:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13200:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13201:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13202:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13203:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13204:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13205:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13206:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd155;
        end
        13207:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        13208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13213:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd161;
        end
        13214:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13215:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13216:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd212;
        end
        13217:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd29;
        end
        13218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13220:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        13221:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13222:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13223:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13224:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13225:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13226:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13227:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13228:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        13229:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        13230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13242:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        13243:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13244:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13245:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13246:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13247:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13248:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13249:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13250:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        13251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13255:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd82;
        end
        13256:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13257:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13258:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13259:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13260:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13261:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13262:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13263:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd217;
        end
        13264:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd30;
        end
        13265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        13317:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd177;
        end
        13318:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13319:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13320:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13321:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13322:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13323:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13324:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13325:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd122;
        end
        13326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13333:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd130;
        end
        13334:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13335:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13336:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13337:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd198;
        end
        13338:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd17;
        end
        13339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13346:
        begin
            RED=8'd0;
            GRN=8'd122;
            BLU=8'd202;
        end
        13347:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13348:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13349:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13350:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13351:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13352:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13353:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13354:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13355:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13356:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13357:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd107;
        end
        13358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13364:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        13365:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        13366:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13367:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13368:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13369:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13370:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13371:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13372:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13373:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13374:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13375:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd38;
        end
        13376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13379:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd102;
        end
        13380:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13381:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13382:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13383:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13384:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13385:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13386:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13387:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13388:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13389:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13390:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        13391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13394:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        13395:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        13396:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13397:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13398:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13399:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13400:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13401:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13402:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13403:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        13404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13428:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd110;
        end
        13429:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13430:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13431:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13432:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13433:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13434:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13435:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13436:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd185;
        end
        13437:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd7;
        end
        13438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13442:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd62;
        end
        13443:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13444:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13445:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13446:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13447:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13448:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13449:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13450:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd210;
        end
        13451:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd27;
        end
        13452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13454:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd177;
        end
        13455:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13456:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13457:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13458:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13459:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13460:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13461:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13462:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd181;
        end
        13463:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd0;
        end
        13464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13469:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd188;
        end
        13470:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13471:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13472:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd205;
        end
        13473:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd20;
        end
        13474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13476:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        13477:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13478:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13479:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13480:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13481:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13482:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13483:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13484:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        13485:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        13486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13498:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        13499:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13500:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13501:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13502:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13503:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13504:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13505:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13506:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        13507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13511:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd68;
        end
        13512:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13513:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13514:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13515:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13516:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13517:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13518:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13519:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd217;
        end
        13520:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd30;
        end
        13521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13572:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd3;
        end
        13573:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        13574:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13575:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13576:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13577:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13578:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13579:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13580:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13581:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd108;
        end
        13582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13589:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd113;
        end
        13590:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        13591:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13592:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13593:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd176;
        end
        13594:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd9;
        end
        13595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd18;
        end
        13602:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd219;
        end
        13603:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13604:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13605:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13606:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13607:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13608:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13609:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13610:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13611:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13612:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13613:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd122;
        end
        13614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13620:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        13621:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        13622:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13623:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13624:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13625:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13626:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13627:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13628:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13629:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13630:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13631:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd76;
        end
        13632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13635:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd131;
        end
        13636:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13637:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13638:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13639:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13640:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13641:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13642:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13643:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13644:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13645:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13646:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        13647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13650:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        13651:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        13652:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13653:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13654:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13655:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13656:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13657:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13658:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13659:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        13660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13684:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd138;
        end
        13685:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13686:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13687:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13688:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13689:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13690:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13691:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13692:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd185;
        end
        13693:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd7;
        end
        13694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13698:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd46;
        end
        13699:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd232;
        end
        13700:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13701:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13702:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13703:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13704:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13705:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13706:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd225;
        end
        13707:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd41;
        end
        13708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13710:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd163;
        end
        13711:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13712:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13713:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13714:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13715:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13716:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13717:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13718:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd203;
        end
        13719:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd13;
        end
        13720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13725:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd202;
        end
        13726:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13727:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13728:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd188;
        end
        13729:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd0;
        end
        13730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13732:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        13733:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13734:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13735:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13736:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13737:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13738:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13739:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13740:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        13741:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        13742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13754:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        13755:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13756:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13757:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13758:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13759:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13760:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13761:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13762:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        13763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13767:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd68;
        end
        13768:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13769:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13770:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13771:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13772:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13773:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13774:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13775:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd217;
        end
        13776:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd30;
        end
        13777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13828:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd24;
        end
        13829:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd231;
        end
        13830:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13831:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13832:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13833:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13834:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13835:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13836:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13837:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd92;
        end
        13838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13845:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd113;
        end
        13846:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        13847:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13848:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd207;
        end
        13849:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd27;
        end
        13850:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        13851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13857:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd42;
        end
        13858:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd224;
        end
        13859:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13860:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13861:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13862:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13863:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13864:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13865:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13866:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13867:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13868:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13869:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd149;
        end
        13870:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        13871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13876:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        13877:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        13878:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13879:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13880:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13881:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13882:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13884:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13885:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13886:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13887:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd90;
        end
        13888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13891:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd157;
        end
        13892:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13893:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13894:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13895:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13896:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13897:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13898:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13899:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13900:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13901:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13902:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        13903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13906:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        13907:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        13908:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13909:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13910:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13911:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13912:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13913:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13914:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13915:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        13916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd3;
        end
        13940:
        begin
            RED=8'd0;
            GRN=8'd95;
            BLU=8'd167;
        end
        13941:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13942:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13943:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13944:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13945:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13946:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13947:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13948:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd172;
        end
        13949:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd4;
        end
        13950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13954:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd46;
        end
        13955:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd232;
        end
        13956:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13957:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13958:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13959:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13960:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13961:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13962:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        13963:
        begin
            RED=8'd0;
            GRN=8'd59;
            BLU=8'd46;
        end
        13964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13966:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd133;
        end
        13967:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13968:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13969:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13970:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13971:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13972:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13973:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13974:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd210;
        end
        13975:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd23;
        end
        13976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd17;
        end
        13981:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd218;
        end
        13982:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13983:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13984:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd162;
        end
        13985:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        13986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13988:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        13989:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13990:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13991:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13992:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13993:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13994:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13995:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        13996:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        13997:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        13998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        13999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14010:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        14011:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14012:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14013:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14014:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14015:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14016:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14017:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14018:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        14019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14023:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd68;
        end
        14024:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14025:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14026:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14027:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14028:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14029:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14030:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14031:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd217;
        end
        14032:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd30;
        end
        14033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14084:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd66;
        end
        14085:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        14086:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14087:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14088:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14089:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14090:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14091:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14092:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14093:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd72;
        end
        14094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14101:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd113;
        end
        14102:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        14103:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd214;
        end
        14104:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd61;
        end
        14105:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd2;
        end
        14106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14113:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd65;
        end
        14114:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd229;
        end
        14115:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14116:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14117:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14118:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14119:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14120:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14121:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14122:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14123:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14124:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14125:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd176;
        end
        14126:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd5;
        end
        14127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14132:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        14133:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        14134:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14135:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14136:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14137:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14138:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14139:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14140:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14141:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14142:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14143:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd116;
        end
        14144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        14147:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd173;
        end
        14148:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14149:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14150:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14151:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14152:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14153:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14154:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14155:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14156:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14157:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14158:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        14159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14162:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        14163:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        14164:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14165:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14166:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14167:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14168:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14169:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14170:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14171:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        14172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd5;
        end
        14196:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd181;
        end
        14197:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14198:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14199:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14200:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14201:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14202:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14203:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14204:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd155;
        end
        14205:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd1;
        end
        14206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14210:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd28;
        end
        14211:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd232;
        end
        14212:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14213:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14214:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14215:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14216:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14217:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14218:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14219:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd81;
        end
        14220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14222:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd101;
        end
        14223:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14224:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14225:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14226:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14227:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14228:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14229:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14230:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd219;
        end
        14231:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd39;
        end
        14232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14236:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd41;
        end
        14237:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd224;
        end
        14238:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14239:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14240:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd135;
        end
        14241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14244:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        14245:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14246:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14247:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14248:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14249:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14250:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14251:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14252:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        14253:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        14254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14266:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        14267:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14268:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14269:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14270:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14271:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14272:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14273:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14274:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        14275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14279:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd82;
        end
        14280:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14281:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14282:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14283:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14284:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14285:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14286:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14287:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd209;
        end
        14288:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd25;
        end
        14289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14340:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd94;
        end
        14341:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14342:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14343:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14344:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14345:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14347:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14348:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd229;
        end
        14349:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd61;
        end
        14350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14357:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd113;
        end
        14358:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd224;
        end
        14359:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd97;
        end
        14360:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd8;
        end
        14361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14369:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd94;
        end
        14370:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd232;
        end
        14371:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14372:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        14373:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd200;
        end
        14374:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14375:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14376:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14377:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14378:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14379:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14380:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14381:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd189;
        end
        14382:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd11;
        end
        14383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14388:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        14389:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        14390:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14391:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14393:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14394:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14396:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14397:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14398:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14399:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd147;
        end
        14400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14402:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd11;
        end
        14403:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd194;
        end
        14404:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14405:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14406:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14407:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14408:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14409:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14410:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14411:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14412:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14413:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14414:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        14415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14418:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        14419:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        14420:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14421:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14422:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14423:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14424:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14425:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14426:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14427:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        14428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14451:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd8;
        end
        14452:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd193;
        end
        14453:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14454:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14455:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14456:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14457:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14458:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14459:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14460:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd153;
        end
        14461:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        14462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14466:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd25;
        end
        14467:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd232;
        end
        14468:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14469:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14470:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14471:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14472:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14473:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14474:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14475:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd98;
        end
        14476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14478:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd85;
        end
        14479:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14480:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14481:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14482:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14483:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14484:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14485:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14486:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd226;
        end
        14487:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd49;
        end
        14488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14492:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd64;
        end
        14493:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd229;
        end
        14494:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14495:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14496:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd118;
        end
        14497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14500:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        14501:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14502:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14503:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14504:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14505:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14506:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14507:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14508:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        14509:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        14510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14522:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        14523:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14524:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14525:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14526:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14527:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14528:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14529:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14530:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        14531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14535:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd96;
        end
        14536:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14537:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14538:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14539:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14540:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14541:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14542:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14543:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd201;
        end
        14544:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd18;
        end
        14545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14596:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd115;
        end
        14597:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14598:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14599:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14600:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14601:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14603:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14604:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        14605:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd59;
        end
        14606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14613:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd48;
        end
        14614:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd82;
        end
        14615:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd20;
        end
        14616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14625:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd113;
        end
        14626:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        14627:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14628:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        14629:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd151;
        end
        14630:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14631:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14632:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14633:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14634:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14635:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14636:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14637:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd207;
        end
        14638:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd18;
        end
        14639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14644:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        14645:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        14646:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14647:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14648:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14649:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14650:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14652:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14653:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14654:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14655:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd178;
        end
        14656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14658:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        14659:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd215;
        end
        14660:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14661:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14662:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14663:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14664:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14665:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14666:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14667:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14668:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14669:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14670:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        14671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14674:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        14675:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        14676:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14677:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14678:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14679:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14680:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14681:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14682:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14683:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        14684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14707:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd12;
        end
        14708:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd214;
        end
        14709:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14710:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14711:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14712:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14713:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14714:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14715:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14716:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd153;
        end
        14717:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        14718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14722:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd25;
        end
        14723:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd232;
        end
        14724:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14725:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14726:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14727:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14728:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14729:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14730:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14731:
        begin
            RED=8'd0;
            GRN=8'd97;
            BLU=8'd112;
        end
        14732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14734:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd61;
        end
        14735:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14736:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14737:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14738:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14739:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14740:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14741:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14742:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        14743:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd72;
        end
        14744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14748:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd77;
        end
        14749:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd231;
        end
        14750:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14751:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        14752:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd89;
        end
        14753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14756:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        14757:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14758:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14759:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14760:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14761:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14762:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14763:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14764:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        14765:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        14766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14778:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        14779:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14780:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14781:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14782:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14783:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14784:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14785:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14786:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        14787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14791:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd109;
        end
        14792:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14793:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14794:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14795:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14796:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14797:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14798:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14799:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd193;
        end
        14800:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd11;
        end
        14801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14852:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd141;
        end
        14853:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14854:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14855:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14856:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14857:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14859:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14860:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd225;
        end
        14861:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd53;
        end
        14862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14869:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd8;
        end
        14870:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd9;
        end
        14871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14881:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd136;
        end
        14882:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14884:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd229;
        end
        14885:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd90;
        end
        14886:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd232;
        end
        14887:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14888:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14889:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14890:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14891:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14892:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14893:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd225;
        end
        14894:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd26;
        end
        14895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14900:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        14901:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        14902:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14903:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14904:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14905:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14906:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14908:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14909:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14910:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14911:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd197;
        end
        14912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14914:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd22;
        end
        14915:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd228;
        end
        14916:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14917:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14918:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14919:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14920:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14921:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14922:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14923:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14924:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14925:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14926:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        14927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14930:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        14931:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        14932:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14933:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14934:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14935:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14936:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14937:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14938:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14939:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        14940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14963:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd14;
        end
        14964:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd228;
        end
        14965:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14966:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14967:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14968:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14969:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14970:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14971:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14972:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd145;
        end
        14973:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd0;
        end
        14974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14978:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd22;
        end
        14979:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd226;
        end
        14980:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14981:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14982:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14983:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14984:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14985:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14986:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14987:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd133;
        end
        14988:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        14989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        14990:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd41;
        end
        14991:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        14992:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14993:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14994:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14995:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14996:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14997:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14998:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        14999:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd101;
        end
        15000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15004:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd104;
        end
        15005:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        15006:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15007:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        15008:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd61;
        end
        15009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15012:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        15013:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15014:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15015:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15016:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15017:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15018:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15019:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15020:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        15021:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        15022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15034:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        15035:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15036:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15037:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15038:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15039:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15040:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15041:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15042:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        15043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15047:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd135;
        end
        15048:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15049:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15050:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15051:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15052:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15053:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15054:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15055:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd166;
        end
        15056:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd3;
        end
        15057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15108:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd162;
        end
        15109:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15110:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15113:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15114:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15115:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15116:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd224;
        end
        15117:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd49;
        end
        15118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15137:
        begin
            RED=8'd0;
            GRN=8'd94;
            BLU=8'd163;
        end
        15138:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15139:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15140:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd221;
        end
        15141:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd49;
        end
        15142:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd228;
        end
        15143:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15144:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15145:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15146:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15147:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15148:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15149:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15150:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd49;
        end
        15151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15156:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        15157:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        15158:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15159:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15161:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15162:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15164:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15165:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15166:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15167:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd218;
        end
        15168:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd0;
        end
        15169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15170:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd44;
        end
        15171:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd232;
        end
        15172:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15173:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15174:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15175:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15176:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15177:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15178:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15179:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15180:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15181:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15182:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        15183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15186:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        15187:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        15188:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15189:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15190:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15191:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15192:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15193:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15194:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15195:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        15196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15219:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd27;
        end
        15220:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd232;
        end
        15221:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15222:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15223:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15224:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15225:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15226:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15227:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15228:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd140;
        end
        15229:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        15230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15234:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd21;
        end
        15235:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd222;
        end
        15236:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15237:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15238:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15239:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15240:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15241:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15242:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15243:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd144;
        end
        15244:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        15245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15246:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd22;
        end
        15247:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd226;
        end
        15248:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15249:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15250:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15251:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15252:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15253:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15254:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15255:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd121;
        end
        15256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15260:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd135;
        end
        15261:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15262:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15263:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd229;
        end
        15264:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd35;
        end
        15265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15268:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        15269:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15270:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15271:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15272:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15273:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15274:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15275:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15276:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        15277:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        15278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15290:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        15291:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15292:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15293:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15294:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15295:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15296:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15297:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15298:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        15299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15303:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd173;
        end
        15304:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15305:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15306:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15307:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15308:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15309:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15310:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15311:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd134;
        end
        15312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15364:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd175;
        end
        15365:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15366:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15367:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15368:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15369:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15370:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15371:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15372:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd222;
        end
        15373:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd44;
        end
        15374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd7;
        end
        15393:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd186;
        end
        15394:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15396:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd208;
        end
        15397:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd31;
        end
        15398:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd218;
        end
        15399:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15400:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15401:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15402:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15403:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15404:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15405:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15406:
        begin
            RED=8'd0;
            GRN=8'd73;
            BLU=8'd74;
        end
        15407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15412:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        15413:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        15414:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15415:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15417:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15418:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15420:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15421:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15422:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15423:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd230;
        end
        15424:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd17;
        end
        15425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15426:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd76;
        end
        15427:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15428:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15429:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15430:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15431:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15432:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15433:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15434:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15435:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15436:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15437:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15438:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        15439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15442:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        15443:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        15444:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15445:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15446:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15447:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15448:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15449:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15450:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15451:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        15452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15475:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd37;
        end
        15476:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd232;
        end
        15477:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15478:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15479:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15480:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15481:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15482:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15483:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15484:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd140;
        end
        15485:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        15486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15490:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd21;
        end
        15491:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd222;
        end
        15492:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15493:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15494:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15495:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15496:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15497:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15498:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15499:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd153;
        end
        15500:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd1;
        end
        15501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15502:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd10;
        end
        15503:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd215;
        end
        15504:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15505:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15506:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15507:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15508:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15509:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15510:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15511:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd140;
        end
        15512:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        15513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15516:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd155;
        end
        15517:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15518:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15519:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd228;
        end
        15520:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd11;
        end
        15521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15524:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        15525:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15526:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15527:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15528:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15529:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15530:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15531:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15532:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        15533:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        15534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15546:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        15547:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15548:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15549:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15550:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15551:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15552:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15553:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15554:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        15555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd16;
        end
        15559:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd209;
        end
        15560:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15561:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15562:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15563:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15564:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15565:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15566:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        15567:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd91;
        end
        15568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15620:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd188;
        end
        15621:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15622:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15623:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15624:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15625:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15626:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15627:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15628:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd220;
        end
        15629:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd39;
        end
        15630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15648:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd21;
        end
        15649:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd205;
        end
        15650:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15652:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd189;
        end
        15653:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd21;
        end
        15654:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd205;
        end
        15655:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15656:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15657:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15658:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15659:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15660:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15661:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15662:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd94;
        end
        15663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15668:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        15669:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        15670:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15671:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15673:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15674:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15676:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15677:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15678:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15679:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        15680:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd44;
        end
        15681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15682:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd102;
        end
        15683:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15684:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15685:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15686:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15687:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15688:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15689:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15690:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15691:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15692:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15693:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15694:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        15695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15698:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        15699:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        15700:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15701:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15702:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15703:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15704:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15705:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15706:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15707:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd66;
        end
        15708:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15709:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15710:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15711:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15712:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15713:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15714:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd18;
        end
        15715:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        15716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15731:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd43;
        end
        15732:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        15733:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15734:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15735:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15736:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15737:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15738:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15739:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15740:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd140;
        end
        15741:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        15742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15746:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd20;
        end
        15747:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd218;
        end
        15748:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15749:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15750:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15751:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15752:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15753:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15754:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15755:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd169;
        end
        15756:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd2;
        end
        15757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15758:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd7;
        end
        15759:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd198;
        end
        15760:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15761:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15762:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15763:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15764:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15765:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15766:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15767:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd162;
        end
        15768:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd2;
        end
        15769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd3;
        end
        15772:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd173;
        end
        15773:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15774:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15775:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd217;
        end
        15776:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd0;
        end
        15777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15780:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        15781:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15782:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15783:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15784:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15785:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15786:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15787:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15788:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        15789:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd50;
        end
        15790:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15791:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15792:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15793:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15794:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15795:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd20;
        end
        15796:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd15;
        end
        15797:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        15798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15802:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        15803:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15804:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15805:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15806:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15807:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15808:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15809:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15810:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        15811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15814:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd69;
        end
        15815:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        15816:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15817:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15818:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15819:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15820:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15821:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15822:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        15823:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd36;
        end
        15824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        15876:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd198;
        end
        15877:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15878:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15879:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15880:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15881:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15882:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15884:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd220;
        end
        15885:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd39;
        end
        15886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15904:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd31;
        end
        15905:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd218;
        end
        15906:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15908:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd159;
        end
        15909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd12;
        end
        15910:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd194;
        end
        15911:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15912:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15913:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15914:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15915:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15916:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15917:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15918:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd122;
        end
        15919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15924:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        15925:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        15926:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15927:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15928:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15929:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15930:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15932:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15933:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15934:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15935:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        15936:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd61;
        end
        15937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15938:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd125;
        end
        15939:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15940:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15941:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15942:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15943:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15944:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15945:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15946:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15947:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15948:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15949:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15950:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        15951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15954:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        15955:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        15956:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15957:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15958:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15959:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15960:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15961:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15962:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15963:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd128;
        end
        15964:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        15965:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        15966:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        15967:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        15968:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        15969:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        15970:
        begin
            RED=8'd0;
            GRN=8'd73;
            BLU=8'd99;
        end
        15971:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd12;
        end
        15972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15987:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd58;
        end
        15988:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15989:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15990:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15991:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15992:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15993:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15994:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15995:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        15996:
        begin
            RED=8'd0;
            GRN=8'd116;
            BLU=8'd136;
        end
        15997:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        15998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        15999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16002:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        16003:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        16004:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16005:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16006:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16007:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16008:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16009:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16010:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16011:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd183;
        end
        16012:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd3;
        end
        16013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        16015:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd172;
        end
        16016:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16017:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16018:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16019:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16020:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16021:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16022:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16023:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd180;
        end
        16024:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd6;
        end
        16025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16027:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd13;
        end
        16028:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd194;
        end
        16029:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16030:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16031:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd191;
        end
        16032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16036:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        16037:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16038:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16039:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16040:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16041:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16042:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16043:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16044:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd222;
        end
        16045:
        begin
            RED=8'd0;
            GRN=8'd94;
            BLU=8'd121;
        end
        16046:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        16047:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        16048:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        16049:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        16050:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        16051:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        16052:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd89;
        end
        16053:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd7;
        end
        16054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16058:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        16059:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16060:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16061:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16062:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16063:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16064:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16065:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16066:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        16067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16069:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd17;
        end
        16070:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd153;
        end
        16071:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        16072:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16073:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16074:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16075:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16076:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16077:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16078:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd194;
        end
        16079:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd0;
        end
        16080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd16;
        end
        16132:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd205;
        end
        16133:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16134:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16135:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16136:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16137:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16138:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16139:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16140:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd219;
        end
        16141:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd37;
        end
        16142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16160:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd41;
        end
        16161:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd226;
        end
        16162:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16164:
        begin
            RED=8'd0;
            GRN=8'd116;
            BLU=8'd129;
        end
        16165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16166:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd176;
        end
        16167:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16168:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16169:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16170:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16171:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16172:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16173:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16174:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd150;
        end
        16175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16180:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        16181:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        16182:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16183:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16185:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16186:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16188:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16189:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16190:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16191:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16192:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd89;
        end
        16193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16194:
        begin
            RED=8'd0;
            GRN=8'd79;
            BLU=8'd148;
        end
        16195:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16196:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16197:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16198:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16199:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16200:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16201:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16202:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16203:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16204:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16205:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16206:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        16207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16210:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        16211:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        16212:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16213:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16214:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16215:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16216:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16217:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16218:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16219:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16220:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16221:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16222:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16223:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16224:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16225:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16226:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd222;
        end
        16227:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd41;
        end
        16228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16243:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd69;
        end
        16244:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16245:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16246:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16247:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16248:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16249:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16250:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16251:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16252:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        16253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16258:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        16259:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        16260:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16261:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16262:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16263:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16264:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16265:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16266:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16267:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd193;
        end
        16268:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd5;
        end
        16269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16271:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd146;
        end
        16272:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16273:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16274:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16275:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16276:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16277:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16278:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16279:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd200;
        end
        16280:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd12;
        end
        16281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16283:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd26;
        end
        16284:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd210;
        end
        16285:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16286:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16287:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd161;
        end
        16288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16292:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        16293:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16294:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16295:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16296:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16297:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16298:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16299:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16300:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16301:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16302:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16303:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16304:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16305:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16306:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16307:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16308:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd207;
        end
        16309:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd22;
        end
        16310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16314:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        16315:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16316:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16317:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16318:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16319:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16320:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16321:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16322:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd164;
        end
        16323:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd11;
        end
        16324:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        16325:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd91;
        end
        16326:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd221;
        end
        16327:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16328:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16329:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16330:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16331:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16332:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16333:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        16334:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd121;
        end
        16335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16387:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd25;
        end
        16388:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd211;
        end
        16389:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16390:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16391:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16393:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16394:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16396:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        16397:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        16398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16416:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd66;
        end
        16417:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        16418:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16420:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd114;
        end
        16421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16422:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd162;
        end
        16423:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16424:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16425:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16426:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16427:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16428:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16429:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16430:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd168;
        end
        16431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16436:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        16437:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        16438:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16439:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16441:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16442:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16443:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16444:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16445:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16446:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16447:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16448:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd120;
        end
        16449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16450:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd177;
        end
        16451:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16452:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16453:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd230;
        end
        16454:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        16455:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16456:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16457:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16458:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16459:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16460:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16461:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16462:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        16463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16466:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        16467:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        16468:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16469:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16470:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16471:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16472:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16473:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16474:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16475:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16476:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16477:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16478:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16479:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16480:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16481:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16482:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd222;
        end
        16483:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd41;
        end
        16484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16499:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd69;
        end
        16500:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16501:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16502:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16503:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16504:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16505:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16506:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16507:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16508:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        16509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16514:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        16515:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        16516:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16517:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16518:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16519:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16520:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16521:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16522:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16523:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd193;
        end
        16524:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd5;
        end
        16525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16527:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd131;
        end
        16528:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16529:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16530:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16531:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16532:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16533:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16534:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16535:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd213;
        end
        16536:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd15;
        end
        16537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16539:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd36;
        end
        16540:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        16541:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16542:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16543:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd129;
        end
        16544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16548:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        16549:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16550:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16551:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16552:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16553:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16554:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16555:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16556:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16557:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16558:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16559:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16560:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16561:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16562:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16563:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16564:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd207;
        end
        16565:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd22;
        end
        16566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16570:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        16571:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16572:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16573:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16574:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16575:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16576:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16577:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16578:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd177;
        end
        16579:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd76;
        end
        16580:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd124;
        end
        16581:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd221;
        end
        16582:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16583:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16584:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16585:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16586:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16587:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16588:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16589:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd210;
        end
        16590:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd37;
        end
        16591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16643:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd34;
        end
        16644:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd216;
        end
        16645:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16646:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16647:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16648:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16649:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16650:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16652:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        16653:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        16654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16655:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd2;
        end
        16656:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16657:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16658:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16659:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16660:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16661:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16662:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16663:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16664:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16665:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16666:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        16667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16672:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd95;
        end
        16673:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16674:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16676:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd87;
        end
        16677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16678:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd134;
        end
        16679:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16680:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16681:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16682:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16683:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16684:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16685:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16686:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd195;
        end
        16687:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        16688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16692:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        16693:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        16694:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16695:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16696:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd229;
        end
        16697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16698:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16699:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16700:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16701:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16702:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16703:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16704:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd150;
        end
        16705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16706:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd203;
        end
        16707:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16708:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16709:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd217;
        end
        16710:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd231;
        end
        16711:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16712:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16713:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16714:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16715:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16716:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16717:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16718:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        16719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16722:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        16723:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        16724:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16725:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16726:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16727:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16728:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16729:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16730:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16731:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16732:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16733:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16734:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16735:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16736:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16737:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16738:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd222;
        end
        16739:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd41;
        end
        16740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16755:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd70;
        end
        16756:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16757:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16758:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16759:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16760:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16761:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16762:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16763:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16764:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        16765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16770:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        16771:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        16772:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16773:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16774:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16775:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16776:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16777:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16778:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16779:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd194;
        end
        16780:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd5;
        end
        16781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16783:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd105;
        end
        16784:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16785:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16786:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16787:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16788:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16789:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16790:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16791:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16792:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd22;
        end
        16793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16795:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd43;
        end
        16796:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd232;
        end
        16797:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16798:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16799:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd116;
        end
        16800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16804:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        16805:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16806:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16807:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16808:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16809:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16810:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16811:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16812:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16813:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16814:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16815:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16816:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16817:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16818:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16819:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16820:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd207;
        end
        16821:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd22;
        end
        16822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16826:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        16827:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16828:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16829:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16830:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16831:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16832:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16833:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16834:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16835:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16836:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16837:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16838:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16839:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16840:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16841:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16842:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16843:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16844:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd230;
        end
        16845:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd126;
        end
        16846:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd0;
        end
        16847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16899:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd34;
        end
        16900:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd216;
        end
        16901:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16902:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16903:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16904:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16905:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16906:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16908:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        16909:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        16910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16911:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd33;
        end
        16912:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16913:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16914:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16915:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16916:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16917:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16918:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16919:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16920:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16921:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16922:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd52;
        end
        16923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        16924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16928:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd123;
        end
        16929:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16930:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16932:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd57;
        end
        16933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16934:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd104;
        end
        16935:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        16936:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16937:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16938:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16939:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16940:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16941:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16942:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd222;
        end
        16943:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd0;
        end
        16944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16948:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        16949:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        16950:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16951:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16952:
        begin
            RED=8'd0;
            GRN=8'd122;
            BLU=8'd174;
        end
        16953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16954:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16955:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16956:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16957:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16958:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16959:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16960:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd164;
        end
        16961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16962:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd216;
        end
        16963:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16964:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16965:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd184;
        end
        16966:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        16967:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16968:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16969:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16970:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16971:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16972:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16973:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16974:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        16975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16978:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        16979:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        16980:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16981:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16982:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16983:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16984:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16985:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16986:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16987:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16988:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16989:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16990:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16991:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16992:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16993:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        16994:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd222;
        end
        16995:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd41;
        end
        16996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        16999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17011:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd84;
        end
        17012:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17013:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17014:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17015:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17016:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17017:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17018:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17019:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17020:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        17021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17026:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        17027:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        17028:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17029:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17030:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17031:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17032:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17033:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17034:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17035:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd207;
        end
        17036:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd6;
        end
        17037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17039:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd91;
        end
        17040:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17041:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17042:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17043:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17044:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17045:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17046:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17047:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17048:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd58;
        end
        17049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17051:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd79;
        end
        17052:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17053:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17054:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17055:
        begin
            RED=8'd0;
            GRN=8'd82;
            BLU=8'd89;
        end
        17056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17060:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        17061:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17062:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17063:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17064:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17065:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17066:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17067:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17068:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17069:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17070:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17071:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17072:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17073:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17074:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17075:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17076:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd207;
        end
        17077:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd22;
        end
        17078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17082:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        17083:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17084:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17085:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17086:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17087:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17088:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17089:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17090:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17091:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17092:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17093:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17094:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17095:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17096:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17097:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17098:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17099:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17100:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd193;
        end
        17101:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd14;
        end
        17102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17155:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd43;
        end
        17156:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd222;
        end
        17157:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17158:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17159:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17161:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17162:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17164:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        17165:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        17166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        17167:
        begin
            RED=8'd0;
            GRN=8'd90;
            BLU=8'd161;
        end
        17168:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17169:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17170:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17171:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17172:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17173:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17174:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17175:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17176:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17177:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17178:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd227;
        end
        17179:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd2;
        end
        17180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17184:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd136;
        end
        17185:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17186:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd224;
        end
        17188:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd31;
        end
        17189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17190:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd83;
        end
        17191:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd232;
        end
        17192:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17193:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17194:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17195:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17196:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17197:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17198:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd224;
        end
        17199:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd18;
        end
        17200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17204:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        17205:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        17206:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17207:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17208:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd137;
        end
        17209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17210:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17211:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17212:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17213:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17214:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17215:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17216:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd190;
        end
        17217:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd31;
        end
        17218:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd222;
        end
        17219:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17220:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17221:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd152;
        end
        17222:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        17223:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17224:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17225:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17226:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17227:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17228:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17229:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17230:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        17231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17234:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        17235:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        17236:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17237:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17238:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17239:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17240:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17241:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17242:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17243:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17244:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17245:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17246:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17247:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17248:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17249:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17250:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd222;
        end
        17251:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd41;
        end
        17252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17267:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd84;
        end
        17268:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17269:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17270:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17271:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17272:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17273:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17274:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17275:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17276:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        17277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17282:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        17283:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        17284:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17285:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17286:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17287:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17288:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17289:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17290:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17291:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd207;
        end
        17292:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd6;
        end
        17293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17295:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd53;
        end
        17296:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd232;
        end
        17297:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17298:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17299:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17300:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17301:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17302:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17303:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17304:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd74;
        end
        17305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17307:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd109;
        end
        17308:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17309:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17310:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17311:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd57;
        end
        17312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17316:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        17317:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17318:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17319:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17320:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17321:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17322:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17323:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17324:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17325:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17326:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17327:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17328:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17329:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17330:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17331:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17332:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd207;
        end
        17333:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd22;
        end
        17334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17338:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        17339:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17340:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17341:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17342:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17343:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17344:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17345:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17347:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17348:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17349:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17350:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17351:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17352:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17353:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17354:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17355:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd206;
        end
        17356:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd30;
        end
        17357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17411:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd43;
        end
        17412:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd222;
        end
        17413:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17414:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17415:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17417:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17418:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17420:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        17421:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        17422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        17423:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd165;
        end
        17424:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17425:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17426:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17427:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17428:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17429:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17430:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17431:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17432:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17433:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17434:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17435:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        17436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17440:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd171;
        end
        17441:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17442:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17443:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd216;
        end
        17444:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd25;
        end
        17445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17446:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd61;
        end
        17447:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd228;
        end
        17448:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17449:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17450:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17451:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17452:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17453:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17454:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd227;
        end
        17455:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd45;
        end
        17456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17460:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        17461:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        17462:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17463:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17464:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd123;
        end
        17465:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17466:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17467:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17468:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17469:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17470:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17471:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17472:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd205;
        end
        17473:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd75;
        end
        17474:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd226;
        end
        17475:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17476:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17477:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd132;
        end
        17478:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        17479:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17480:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17481:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17482:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17483:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17484:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17485:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17486:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        17487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17490:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        17491:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        17492:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17493:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17494:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17495:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17496:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17497:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17498:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17499:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17500:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17501:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17502:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17503:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17504:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17505:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17506:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd222;
        end
        17507:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd41;
        end
        17508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17523:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd84;
        end
        17524:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17525:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17526:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17527:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17528:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17529:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17530:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17531:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17532:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        17533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17538:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        17539:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        17540:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17541:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17542:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17543:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17544:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17545:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17546:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17547:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd207;
        end
        17548:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd6;
        end
        17549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17551:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd39;
        end
        17552:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd220;
        end
        17553:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17554:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17555:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17556:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17557:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17558:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17559:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17560:
        begin
            RED=8'd0;
            GRN=8'd94;
            BLU=8'd100;
        end
        17561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17563:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd134;
        end
        17564:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17565:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17566:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd224;
        end
        17567:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd33;
        end
        17568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17572:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        17573:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17574:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17575:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17576:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17577:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17578:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17579:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17580:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17581:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17582:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17583:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17584:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17585:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17586:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17587:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17588:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd207;
        end
        17589:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd22;
        end
        17590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17594:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        17595:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17596:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17597:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17598:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17599:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17600:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17601:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17603:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17604:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17605:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17606:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17607:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17608:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17609:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17610:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd185;
        end
        17611:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd31;
        end
        17612:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        17613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17667:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd43;
        end
        17668:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd222;
        end
        17669:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17670:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17671:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17673:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17674:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17676:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        17677:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        17678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        17679:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd165;
        end
        17680:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17681:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17682:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17683:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17684:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17685:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17686:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17687:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17688:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17689:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17690:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17691:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        17692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        17696:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd199;
        end
        17697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17698:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17699:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd199;
        end
        17700:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd16;
        end
        17701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17702:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd48;
        end
        17703:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd226;
        end
        17704:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17705:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17706:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17707:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17708:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17709:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17710:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        17711:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd69;
        end
        17712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17716:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        17717:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        17718:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17719:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17720:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd98;
        end
        17721:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17722:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17723:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17724:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17725:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17726:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17727:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17728:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd213;
        end
        17729:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd105;
        end
        17730:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd231;
        end
        17731:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17732:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        17733:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd108;
        end
        17734:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        17735:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17736:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17737:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17738:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17739:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17740:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17741:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17742:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        17743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17746:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        17747:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        17748:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17749:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17750:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17751:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17752:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17753:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17754:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17755:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd88;
        end
        17756:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17757:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17758:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17759:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17760:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17761:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17762:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd42;
        end
        17763:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd8;
        end
        17764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17779:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd84;
        end
        17780:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17781:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17782:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17783:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17784:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17785:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17786:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17787:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17788:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        17789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17794:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        17795:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        17796:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17797:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17798:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17799:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17800:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17801:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17802:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17803:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd207;
        end
        17804:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd6;
        end
        17805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17807:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd30;
        end
        17808:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd214;
        end
        17809:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17810:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17811:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17812:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17813:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17814:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17815:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17816:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd113;
        end
        17817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17819:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd154;
        end
        17820:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17821:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17822:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd216;
        end
        17823:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd26;
        end
        17824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17828:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        17829:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17830:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17831:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17832:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17833:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17834:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17835:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17836:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd221;
        end
        17837:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd73;
        end
        17838:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17839:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17840:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17841:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17842:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17843:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd44;
        end
        17844:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd39;
        end
        17845:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd4;
        end
        17846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17850:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        17851:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17852:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17853:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17854:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17855:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17856:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17857:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17859:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17860:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17861:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17862:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17863:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17864:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17865:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17866:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd222;
        end
        17867:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd111;
        end
        17868:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        17869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17923:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd43;
        end
        17924:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd222;
        end
        17925:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17926:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17927:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17928:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17929:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17930:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17932:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        17933:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        17934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        17935:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd165;
        end
        17936:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17937:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17938:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17939:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17940:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17941:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17942:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17943:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17944:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17945:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17946:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17947:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        17948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        17952:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd224;
        end
        17953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17954:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17955:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd177;
        end
        17956:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd4;
        end
        17957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17958:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd25;
        end
        17959:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd222;
        end
        17960:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17961:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17962:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17963:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17964:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17965:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17966:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        17967:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd83;
        end
        17968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        17972:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        17973:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        17974:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17975:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17976:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd69;
        end
        17977:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd232;
        end
        17978:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17979:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17980:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17981:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17982:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17983:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17984:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd223;
        end
        17985:
        begin
            RED=8'd0;
            GRN=8'd94;
            BLU=8'd139;
        end
        17986:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        17987:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17988:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd229;
        end
        17989:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd82;
        end
        17990:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        17991:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17992:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17993:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17994:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17995:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17996:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17997:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        17998:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        17999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18002:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        18003:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        18004:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18005:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18006:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18007:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18008:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18009:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18010:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18011:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        18012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18035:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd84;
        end
        18036:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18037:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18038:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18039:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18040:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18041:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18042:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18043:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18044:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        18045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18050:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        18051:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        18052:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18053:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18054:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18055:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18056:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18057:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18058:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18059:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd207;
        end
        18060:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd6;
        end
        18061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18063:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd17;
        end
        18064:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd202;
        end
        18065:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18066:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18067:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18068:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18069:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18070:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18071:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18072:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd144;
        end
        18073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        18075:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd181;
        end
        18076:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18077:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18078:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd200;
        end
        18079:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd17;
        end
        18080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18084:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        18085:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18086:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18087:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18088:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18089:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18090:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18091:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18092:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        18093:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        18094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18106:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        18107:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18108:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18109:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18110:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18113:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18114:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd182;
        end
        18115:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd63;
        end
        18116:
        begin
            RED=8'd0;
            GRN=8'd95;
            BLU=8'd158;
        end
        18117:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18118:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18119:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18120:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18121:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18122:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18123:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd206;
        end
        18124:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd55;
        end
        18125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18179:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd43;
        end
        18180:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd222;
        end
        18181:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18182:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18183:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18185:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18186:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18188:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        18189:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        18190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        18191:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd165;
        end
        18192:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18193:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18194:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18195:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18196:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18197:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18198:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18199:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18200:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18201:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18202:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18203:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        18204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18207:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd26;
        end
        18208:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd232;
        end
        18209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18210:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18211:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd162;
        end
        18212:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd0;
        end
        18213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd6;
        end
        18215:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd210;
        end
        18216:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18217:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18218:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18219:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18220:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18221:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18222:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18223:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd111;
        end
        18224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18228:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        18229:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        18230:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18231:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18232:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd45;
        end
        18233:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd225;
        end
        18234:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18235:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18236:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18237:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18238:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18239:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18240:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        18241:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd203;
        end
        18242:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        18243:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18244:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd228;
        end
        18245:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd65;
        end
        18246:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        18247:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18248:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18249:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18250:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18251:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18252:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18253:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18254:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        18255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18258:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        18259:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        18260:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18261:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18262:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18263:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18264:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18265:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18266:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18267:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        18268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18291:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd84;
        end
        18292:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18293:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18294:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18295:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18296:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18297:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18298:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18299:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18300:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        18301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18306:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        18307:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        18308:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18309:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18310:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18311:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18312:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18313:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18314:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18315:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd207;
        end
        18316:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd6;
        end
        18317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        18320:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd191;
        end
        18321:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18322:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18323:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18324:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18325:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18326:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18327:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18328:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd164;
        end
        18329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18330:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        18331:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd209;
        end
        18332:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18333:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18334:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd179;
        end
        18335:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd5;
        end
        18336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18340:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        18341:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18342:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18343:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18344:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18345:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18347:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18348:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        18349:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        18350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18362:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        18363:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18364:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18365:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18366:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18367:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18368:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18369:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18370:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        18371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18372:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd47;
        end
        18373:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd179;
        end
        18374:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18375:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18376:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18377:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18378:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18379:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18380:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd164;
        end
        18381:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd16;
        end
        18382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18435:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd43;
        end
        18436:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd222;
        end
        18437:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18438:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18439:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18441:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18442:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18443:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18444:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        18445:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        18446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        18447:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd165;
        end
        18448:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18449:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18450:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18451:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18452:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18453:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18454:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18455:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18456:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18457:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18458:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18459:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        18460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18463:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd48;
        end
        18464:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18465:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18466:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18467:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd140;
        end
        18468:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        18469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18471:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd197;
        end
        18472:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18473:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18474:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18475:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18476:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18477:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18478:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18479:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd142;
        end
        18480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18484:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        18485:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        18486:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18487:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18488:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd35;
        end
        18489:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd214;
        end
        18490:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18491:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18492:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18493:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18494:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18495:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18496:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18497:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18498:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18499:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18500:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd220;
        end
        18501:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd47;
        end
        18502:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        18503:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18504:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18505:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18506:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18507:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18508:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18509:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18510:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        18511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18514:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        18515:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        18516:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18517:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18518:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18519:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18520:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18521:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18522:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18523:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        18524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18547:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd75;
        end
        18548:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18549:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18550:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18551:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18552:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18553:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18554:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18555:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18556:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        18557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18562:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        18563:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        18564:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18565:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18566:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18567:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18568:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18569:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18570:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18571:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd207;
        end
        18572:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd6;
        end
        18573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18576:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd172;
        end
        18577:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18578:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18579:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18580:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18581:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18582:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18583:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18584:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd186;
        end
        18585:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd0;
        end
        18586:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        18587:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd226;
        end
        18588:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18589:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18590:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd155;
        end
        18591:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd0;
        end
        18592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18596:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        18597:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18598:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18599:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18600:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18601:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18603:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18604:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        18605:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        18606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18618:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        18619:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18620:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18621:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18622:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18623:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18624:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18625:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18626:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        18627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        18629:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd92;
        end
        18630:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd232;
        end
        18631:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18632:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18633:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18634:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18635:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18636:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd223;
        end
        18637:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd86;
        end
        18638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18691:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd39;
        end
        18692:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd219;
        end
        18693:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18694:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18695:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18696:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18698:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18699:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18700:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        18701:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        18702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        18703:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd85;
        end
        18704:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd119;
        end
        18705:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd119;
        end
        18706:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd119;
        end
        18707:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd219;
        end
        18708:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18709:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18710:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18711:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18712:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18713:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18714:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18715:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        18716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18719:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd69;
        end
        18720:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18721:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18722:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18723:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd112;
        end
        18724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18727:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd176;
        end
        18728:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18729:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18730:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18731:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18732:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18733:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18734:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18735:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd162;
        end
        18736:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        18737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18740:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        18741:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        18742:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18743:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18744:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd31;
        end
        18745:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd197;
        end
        18746:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18747:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18748:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18749:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18750:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18751:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18752:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18753:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18754:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18755:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18756:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd200;
        end
        18757:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd38;
        end
        18758:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        18759:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18760:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18761:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18762:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18763:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18764:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18765:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18766:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        18767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18770:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        18771:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        18772:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18773:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18774:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18775:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18776:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18777:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18778:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18779:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        18780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18803:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd69;
        end
        18804:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18805:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18806:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18807:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18808:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18809:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18810:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18811:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18812:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        18813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18818:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        18819:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        18820:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18821:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18822:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18823:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18824:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18825:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18826:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18827:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd200;
        end
        18828:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd5;
        end
        18829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18832:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd145;
        end
        18833:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18834:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18835:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18836:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18837:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18838:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18839:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18840:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd208;
        end
        18841:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd8;
        end
        18842:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd20;
        end
        18843:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd232;
        end
        18844:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18845:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18846:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd136;
        end
        18847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18852:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        18853:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18854:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18855:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18856:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18857:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18859:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18860:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        18861:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        18862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18874:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        18875:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18876:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18877:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18878:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18879:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18880:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18881:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18882:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        18883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18885:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd30;
        end
        18886:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd213;
        end
        18887:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18888:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18889:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18890:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18891:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18892:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18893:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd170;
        end
        18894:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd8;
        end
        18895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18947:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd34;
        end
        18948:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd216;
        end
        18949:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18950:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18951:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18952:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18954:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18955:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18956:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        18957:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        18958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18963:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        18964:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18965:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18966:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18967:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18968:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18969:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18970:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18971:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        18972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18975:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd98;
        end
        18976:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18977:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18978:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        18979:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd83;
        end
        18980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18983:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd153;
        end
        18984:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18985:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18986:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18987:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18988:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18989:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18990:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18991:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd179;
        end
        18992:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd4;
        end
        18993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        18996:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        18997:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        18998:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        18999:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19000:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd26;
        end
        19001:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd171;
        end
        19002:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19003:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19004:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19005:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19006:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19007:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19008:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19009:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19010:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19011:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19012:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd178;
        end
        19013:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        19014:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        19015:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19016:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19017:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19018:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19019:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19020:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19021:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19022:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        19023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19026:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        19027:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        19028:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19029:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19030:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19031:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19032:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19033:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19034:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19035:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        19036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19059:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd69;
        end
        19060:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19061:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19062:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19063:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19064:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19065:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19066:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19067:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19068:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        19069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19074:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        19075:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        19076:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19077:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19078:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19079:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19080:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19081:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19082:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19083:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd193;
        end
        19084:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd5;
        end
        19085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19088:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd123;
        end
        19089:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19090:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19091:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19092:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19093:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19094:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19095:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19096:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd218;
        end
        19097:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd23;
        end
        19098:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd52;
        end
        19099:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19100:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19101:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19102:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd115;
        end
        19103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19108:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        19109:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19110:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19113:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19114:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19115:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19116:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        19117:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        19118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19130:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        19131:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19132:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19133:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19134:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19135:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19136:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19137:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19138:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        19139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd7;
        end
        19142:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd178;
        end
        19143:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19144:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19145:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19146:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19147:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19148:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19149:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        19150:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd36;
        end
        19151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19203:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd31;
        end
        19204:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd214;
        end
        19205:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19206:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19207:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19208:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19210:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19211:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19212:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        19213:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        19214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19219:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        19220:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19221:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19222:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19223:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19224:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19225:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19226:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19227:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        19228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19231:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd129;
        end
        19232:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19233:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19234:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        19235:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd60;
        end
        19236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19239:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd132;
        end
        19240:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19241:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19242:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19243:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19244:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19245:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19246:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19247:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd199;
        end
        19248:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd16;
        end
        19249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19252:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        19253:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        19254:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19255:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19256:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        19257:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd143;
        end
        19258:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19259:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19260:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19261:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19262:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19263:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19264:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19265:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19266:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19267:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19268:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd156;
        end
        19269:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        19270:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        19271:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19272:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19273:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19274:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19275:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19276:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19277:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19278:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        19279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19282:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        19283:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        19284:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19285:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19286:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19287:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19288:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19289:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19290:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19291:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        19292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19315:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd64;
        end
        19316:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19317:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19318:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19319:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19320:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19321:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19322:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19323:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19324:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd126;
        end
        19325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19330:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd18;
        end
        19331:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        19332:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19333:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19334:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19335:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19336:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19337:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19338:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19339:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd188;
        end
        19340:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd4;
        end
        19341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19344:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd102;
        end
        19345:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        19346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19347:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19348:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19349:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19350:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19351:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19352:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd222;
        end
        19353:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd39;
        end
        19354:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd79;
        end
        19355:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19356:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19357:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        19358:
        begin
            RED=8'd0;
            GRN=8'd82;
            BLU=8'd85;
        end
        19359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19364:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        19365:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19366:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19367:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19368:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19369:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19370:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19371:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19372:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        19373:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        19374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19386:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        19387:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19388:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19389:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19390:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19391:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19393:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19394:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        19395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19398:
        begin
            RED=8'd0;
            GRN=8'd79;
            BLU=8'd146;
        end
        19399:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19400:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19401:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19402:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19403:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19404:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19405:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19406:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd77;
        end
        19407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd24;
        end
        19460:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd210;
        end
        19461:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19462:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19463:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19464:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19465:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19466:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19467:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19468:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        19469:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd28;
        end
        19470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19475:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        19476:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19477:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19478:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19479:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19480:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19481:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19482:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19483:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        19484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19487:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd158;
        end
        19488:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19489:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19490:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd224;
        end
        19491:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd47;
        end
        19492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19495:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd104;
        end
        19496:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19497:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19498:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19499:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19500:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19501:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19502:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19503:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd212;
        end
        19504:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd28;
        end
        19505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19508:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        19509:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        19510:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19511:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19512:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        19513:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd121;
        end
        19514:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19515:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19516:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19517:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19518:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19519:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19520:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19521:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19522:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19523:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19524:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd124;
        end
        19525:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        19526:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        19527:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19528:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19529:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19530:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19531:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19532:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19533:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19534:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        19535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19538:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        19539:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        19540:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19541:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19542:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19543:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19544:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19545:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19546:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19547:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        19548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19571:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd50;
        end
        19572:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        19573:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19574:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19575:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19576:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19577:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19578:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19579:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19580:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd129;
        end
        19581:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        19582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19586:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd19;
        end
        19587:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd214;
        end
        19588:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19589:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19590:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19591:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19592:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19593:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19594:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19595:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd179;
        end
        19596:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd3;
        end
        19597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19600:
        begin
            RED=8'd0;
            GRN=8'd33;
            BLU=8'd76;
        end
        19601:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd231;
        end
        19602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19603:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19604:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19605:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19606:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19607:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19608:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd227;
        end
        19609:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd58;
        end
        19610:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd103;
        end
        19611:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19612:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19613:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd227;
        end
        19614:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd58;
        end
        19615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19620:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        19621:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19622:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19623:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19624:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19625:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19626:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19627:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19628:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        19629:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        19630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19642:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        19643:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19644:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19645:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19646:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19647:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19648:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19649:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19650:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        19651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19654:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd116;
        end
        19655:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        19656:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19657:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19658:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19659:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19660:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19661:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19662:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd115;
        end
        19663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd22;
        end
        19716:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd209;
        end
        19717:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19718:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19719:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19720:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19721:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19722:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19723:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19724:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd216;
        end
        19725:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd30;
        end
        19726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19731:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        19732:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19733:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19734:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19735:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19736:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19737:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19738:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19739:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        19740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19743:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd182;
        end
        19744:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19745:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19746:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd217;
        end
        19747:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd25;
        end
        19748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19751:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd89;
        end
        19752:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19753:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19754:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19755:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19756:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19757:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19758:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19759:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd220;
        end
        19760:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd36;
        end
        19761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19764:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        19765:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        19766:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19767:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19768:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        19769:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd104;
        end
        19770:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        19771:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19772:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19773:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19774:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19775:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19776:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19777:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19778:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19779:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19780:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd101;
        end
        19781:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        19782:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        19783:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19784:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19785:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19786:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19787:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19788:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19789:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19790:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        19791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19794:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        19795:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        19796:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19797:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19798:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19799:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19800:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19801:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19802:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19803:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        19804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19827:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd37;
        end
        19828:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd232;
        end
        19829:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19830:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19831:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19832:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19833:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19834:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19835:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19836:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd140;
        end
        19837:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        19838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19842:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd21;
        end
        19843:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd222;
        end
        19844:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19845:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19846:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19847:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19848:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19849:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19850:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19851:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd176;
        end
        19852:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd3;
        end
        19853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19856:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd60;
        end
        19857:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd231;
        end
        19858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19859:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19860:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19861:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19862:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19863:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19864:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd229;
        end
        19865:
        begin
            RED=8'd0;
            GRN=8'd73;
            BLU=8'd71;
        end
        19866:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd124;
        end
        19867:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19868:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19869:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd222;
        end
        19870:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd39;
        end
        19871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19876:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        19877:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19878:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19879:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19880:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19881:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19882:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19884:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        19885:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        19886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19898:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        19899:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19900:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19901:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19902:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19903:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19904:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19905:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19906:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        19907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19910:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd85;
        end
        19911:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        19912:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19913:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19914:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19915:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19916:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19917:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19918:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd147;
        end
        19919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd13;
        end
        19972:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd203;
        end
        19973:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19974:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19975:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19976:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19977:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19978:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19979:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19980:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd220;
        end
        19981:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd39;
        end
        19982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19987:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        19988:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19989:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19990:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19991:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19992:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19993:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19994:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        19995:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        19996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        19998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        19999:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd195;
        end
        20000:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20001:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20002:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd209;
        end
        20003:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd0;
        end
        20004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20007:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd61;
        end
        20008:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        20009:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20010:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20011:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20012:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20013:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20014:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20015:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20016:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd50;
        end
        20017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20020:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        20021:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        20022:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20023:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20024:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        20025:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd75;
        end
        20026:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd231;
        end
        20027:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20028:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20029:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20030:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20031:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20032:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20033:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20034:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20035:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20036:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd85;
        end
        20037:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        20038:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        20039:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20040:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20041:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20042:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20043:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20044:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20045:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20046:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        20047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20050:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        20051:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        20052:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20053:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20054:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20055:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20056:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20057:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20058:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20059:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        20060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20083:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd35;
        end
        20084:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd232;
        end
        20085:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20086:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20087:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20088:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20089:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20090:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20091:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20092:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd140;
        end
        20093:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        20094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20098:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd21;
        end
        20099:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd222;
        end
        20100:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20101:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20102:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20103:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20104:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20105:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20106:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20107:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd161;
        end
        20108:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd2;
        end
        20109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd34;
        end
        20113:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd229;
        end
        20114:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20115:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20116:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20117:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20118:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20119:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20120:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20121:
        begin
            RED=8'd0;
            GRN=8'd94;
            BLU=8'd101;
        end
        20122:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd154;
        end
        20123:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20124:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20125:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd218;
        end
        20126:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd28;
        end
        20127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20132:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        20133:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20134:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20135:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20136:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20137:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20138:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20139:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20140:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        20141:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        20142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20154:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        20155:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20156:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20157:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20158:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20159:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20161:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20162:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        20163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20166:
        begin
            RED=8'd0;
            GRN=8'd33;
            BLU=8'd74;
        end
        20167:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd231;
        end
        20168:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20169:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20170:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20171:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20172:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20173:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20174:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd177;
        end
        20175:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        20176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20228:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd196;
        end
        20229:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20230:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20231:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20232:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20233:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20234:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20235:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20236:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd220;
        end
        20237:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd39;
        end
        20238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20243:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        20244:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20245:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20246:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20247:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20248:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20249:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20250:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20251:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        20252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd23;
        end
        20255:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd209;
        end
        20256:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20257:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20258:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd197;
        end
        20259:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd0;
        end
        20260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20263:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd25;
        end
        20264:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd232;
        end
        20265:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20266:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20267:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20268:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20269:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20270:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20271:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20272:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd85;
        end
        20273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20276:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        20277:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        20278:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20279:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20280:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        20281:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd48;
        end
        20282:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd226;
        end
        20283:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20284:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20285:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20286:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20287:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20288:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20289:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20290:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20291:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20292:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd56;
        end
        20293:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        20294:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        20295:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20296:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20297:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20298:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20299:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20300:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20301:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20302:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        20303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20306:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        20307:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        20308:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20309:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20310:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20311:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20312:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20313:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20314:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20315:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        20316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20339:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd15;
        end
        20340:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd232;
        end
        20341:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20342:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20343:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20344:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20345:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20347:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20348:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd140;
        end
        20349:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        20350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20354:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd21;
        end
        20355:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd222;
        end
        20356:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20357:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20358:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20359:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20360:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20361:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20362:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20363:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd144;
        end
        20364:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        20365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20369:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd227;
        end
        20370:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20371:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20372:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20373:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20374:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20375:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20376:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20377:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd131;
        end
        20378:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd181;
        end
        20379:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20380:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20381:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd209;
        end
        20382:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd0;
        end
        20383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20388:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        20389:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20390:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20391:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20393:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20394:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20396:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        20397:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        20398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20410:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        20411:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20412:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20413:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20414:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20415:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20417:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20418:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        20419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20422:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd62;
        end
        20423:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd229;
        end
        20424:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20425:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20426:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20427:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20428:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20429:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20430:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd204;
        end
        20431:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd0;
        end
        20432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20484:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd183;
        end
        20485:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20486:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20487:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20488:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20489:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20490:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20491:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20492:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd220;
        end
        20493:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd39;
        end
        20494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20499:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        20500:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20501:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20502:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20503:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20504:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20505:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20506:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20507:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        20508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20510:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd42;
        end
        20511:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd221;
        end
        20512:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20513:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20514:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd168;
        end
        20515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20519:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd22;
        end
        20520:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd222;
        end
        20521:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20522:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20523:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20524:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20525:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20526:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20527:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20528:
        begin
            RED=8'd0;
            GRN=8'd90;
            BLU=8'd101;
        end
        20529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20532:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        20533:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        20534:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20535:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20536:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        20537:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd31;
        end
        20538:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd214;
        end
        20539:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20540:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20541:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20542:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20543:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20544:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20545:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20546:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20547:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd223;
        end
        20548:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd30;
        end
        20549:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        20550:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        20551:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20552:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20553:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20554:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20555:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20556:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20557:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20558:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        20559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20562:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        20563:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        20564:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20565:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20566:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20567:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20568:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20569:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20570:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20571:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        20572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20595:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd13;
        end
        20596:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd221;
        end
        20597:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20598:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20599:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20600:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20601:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20603:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20604:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd140;
        end
        20605:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        20606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20610:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd21;
        end
        20611:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd222;
        end
        20612:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20613:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20614:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20615:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20616:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20617:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20618:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20619:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd130;
        end
        20620:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        20621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20625:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd214;
        end
        20626:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20627:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20628:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20629:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20630:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20631:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20632:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20633:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd159;
        end
        20634:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd203;
        end
        20635:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20636:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20637:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd182;
        end
        20638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20644:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        20645:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20646:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20647:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20648:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20649:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20650:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20652:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        20653:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        20654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20666:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        20667:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20668:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20669:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20670:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20671:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20673:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20674:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        20675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20678:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd49;
        end
        20679:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        20680:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20681:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20682:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20683:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20684:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20685:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20686:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd217;
        end
        20687:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd0;
        end
        20688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20740:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd156;
        end
        20741:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20742:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20743:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20744:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20745:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20746:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20747:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20748:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd224;
        end
        20749:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd48;
        end
        20750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20755:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        20756:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20757:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20758:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20759:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20760:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20761:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20762:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20763:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        20764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20766:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd57;
        end
        20767:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd231;
        end
        20768:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20769:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20770:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd158;
        end
        20771:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd48;
        end
        20772:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd48;
        end
        20773:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd48;
        end
        20774:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd48;
        end
        20775:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd61;
        end
        20776:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd213;
        end
        20777:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20778:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20779:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20780:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20781:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20782:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20783:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20784:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd127;
        end
        20785:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        20786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20788:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        20789:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        20790:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20791:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20792:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        20793:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd23;
        end
        20794:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd208;
        end
        20795:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20796:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20797:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20798:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20799:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20800:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20801:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20802:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20803:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd215;
        end
        20804:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd24;
        end
        20805:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        20806:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        20807:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20808:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20809:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20810:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20811:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20812:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20813:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20814:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        20815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20818:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        20819:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        20820:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20821:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20822:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20823:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20824:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20825:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20826:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20827:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        20828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20851:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd9;
        end
        20852:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd198;
        end
        20853:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20854:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20855:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20856:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20857:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20859:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20860:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd152;
        end
        20861:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        20862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20866:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd24;
        end
        20867:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd231;
        end
        20868:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20869:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20870:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20871:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20872:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20873:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20874:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20875:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd117;
        end
        20876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20881:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd187;
        end
        20882:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20884:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20885:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20886:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20887:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20888:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20889:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd202;
        end
        20890:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd214;
        end
        20891:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20892:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20893:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd154;
        end
        20894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20900:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        20901:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20902:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20903:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20904:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20905:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20906:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20908:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        20909:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        20910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20922:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        20923:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20924:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20925:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20926:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20927:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20928:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20929:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20930:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        20931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20934:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd49;
        end
        20935:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        20936:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20937:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20938:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20939:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20940:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20941:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20942:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd220;
        end
        20943:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd17;
        end
        20944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        20996:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd140;
        end
        20997:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20998:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        20999:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21000:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21001:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21002:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21003:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21004:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd224;
        end
        21005:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd49;
        end
        21006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21011:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        21012:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21013:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21014:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21015:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21016:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21017:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21018:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21019:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        21020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21022:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd76;
        end
        21023:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        21024:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21025:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21026:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd220;
        end
        21027:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd203;
        end
        21028:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd203;
        end
        21029:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd203;
        end
        21030:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd203;
        end
        21031:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd205;
        end
        21032:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd229;
        end
        21033:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21034:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21035:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21036:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21037:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21038:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21039:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21040:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd158;
        end
        21041:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd2;
        end
        21042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21044:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        21045:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        21046:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21047:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21048:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        21049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        21050:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd194;
        end
        21051:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21052:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21053:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21054:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21055:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21056:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21057:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21058:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21059:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd198;
        end
        21060:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd15;
        end
        21061:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        21062:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        21063:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21064:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21065:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21066:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21067:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21068:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21069:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21070:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        21071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21074:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        21075:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        21076:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21077:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21078:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21079:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21080:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21081:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21082:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21083:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        21084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd6;
        end
        21108:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd185;
        end
        21109:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21110:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21113:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21114:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21115:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21116:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd153;
        end
        21117:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        21118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21122:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd25;
        end
        21123:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd232;
        end
        21124:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21125:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21126:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21127:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21128:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21129:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21130:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21131:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd103;
        end
        21132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21137:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd171;
        end
        21138:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21139:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21140:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21141:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21142:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21143:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21144:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21145:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd228;
        end
        21146:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd229;
        end
        21147:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21148:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21149:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd138;
        end
        21150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21156:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        21157:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21158:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21159:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21161:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21162:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21164:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        21165:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        21166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21178:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        21179:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21180:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21181:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21182:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21183:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21185:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21186:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        21187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21190:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd49;
        end
        21191:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        21192:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21193:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21194:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21195:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21196:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21197:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21198:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd222;
        end
        21199:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd30;
        end
        21200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21252:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd109;
        end
        21253:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21254:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21255:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21256:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21257:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21258:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21259:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21260:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd227;
        end
        21261:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd56;
        end
        21262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21267:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        21268:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21269:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21270:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21271:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21272:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21273:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21274:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21275:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        21276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21278:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd104;
        end
        21279:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        21280:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21281:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21282:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21283:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21284:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21285:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21286:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21287:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21288:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21289:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21290:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21291:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21292:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21293:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21294:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21295:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21296:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd175;
        end
        21297:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd3;
        end
        21298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21300:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        21301:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        21302:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21303:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21304:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        21305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21306:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd170;
        end
        21307:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21308:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21309:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21310:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21311:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21312:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21313:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21314:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21315:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd176;
        end
        21316:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd3;
        end
        21317:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        21318:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        21319:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21320:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21321:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21322:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21323:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21324:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21325:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21326:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        21327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21330:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        21331:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        21332:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21333:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21334:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21335:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21336:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21337:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21338:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21339:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        21340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        21364:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd172;
        end
        21365:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21366:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21367:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21368:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21369:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21370:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21371:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21372:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd166;
        end
        21373:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd3;
        end
        21374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21378:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd25;
        end
        21379:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd232;
        end
        21380:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21381:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21382:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21383:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21384:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21385:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21386:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21387:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd77;
        end
        21388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21393:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd140;
        end
        21394:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21396:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21397:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21398:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21399:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21400:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21401:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21402:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21403:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21404:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21405:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd108;
        end
        21406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21412:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        21413:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21414:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21415:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21417:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21418:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21420:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        21421:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        21422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21434:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        21435:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21436:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21437:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21438:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21439:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21441:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21442:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        21443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21446:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd49;
        end
        21447:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        21448:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21449:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21450:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21451:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21452:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21453:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21454:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        21455:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd43;
        end
        21456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21508:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd81;
        end
        21509:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21510:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21511:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21512:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21513:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21514:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21515:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21516:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        21517:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd59;
        end
        21518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21523:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        21524:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21525:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21526:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21527:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21528:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21529:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21530:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21531:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        21532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21534:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd132;
        end
        21535:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21536:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21537:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21538:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21539:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21540:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21541:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21542:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21543:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21544:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21545:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21546:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21547:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21548:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21549:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21550:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21551:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21552:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd198;
        end
        21553:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd4;
        end
        21554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21556:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        21557:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        21558:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21559:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21560:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        21561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21562:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd144;
        end
        21563:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21564:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21565:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21566:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21567:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21568:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21569:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21570:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21571:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd161;
        end
        21572:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd0;
        end
        21573:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        21574:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        21575:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21576:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21577:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21578:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21579:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21580:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21581:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21582:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        21583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21586:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        21587:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        21588:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21589:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21590:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21591:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21592:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21593:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21594:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21595:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        21596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        21620:
        begin
            RED=8'd0;
            GRN=8'd82;
            BLU=8'd148;
        end
        21621:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21622:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21623:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21624:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21625:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21626:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21627:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21628:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd171;
        end
        21629:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd4;
        end
        21630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21634:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd39;
        end
        21635:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd232;
        end
        21636:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21637:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21638:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21639:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21640:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21641:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21642:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21643:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd54;
        end
        21644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21649:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd112;
        end
        21650:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21652:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21653:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21654:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21655:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21656:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21657:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21658:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21659:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21660:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21661:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd80;
        end
        21662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21668:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        21669:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21670:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21671:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21673:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21674:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21676:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        21677:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        21678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21690:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        21691:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21692:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21693:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21694:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21695:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21696:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21698:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        21699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21702:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd49;
        end
        21703:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        21704:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21705:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21706:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21707:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21708:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21709:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21710:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd227;
        end
        21711:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd54;
        end
        21712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21764:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd54;
        end
        21765:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21766:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21767:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21768:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21769:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21770:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21771:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21772:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        21773:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd65;
        end
        21774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21779:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        21780:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21781:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21782:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21783:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21784:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21785:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21786:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21787:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        21788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        21790:
        begin
            RED=8'd0;
            GRN=8'd90;
            BLU=8'd159;
        end
        21791:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21792:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21793:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21794:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21795:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21796:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21797:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21798:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21799:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21800:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21801:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21802:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21803:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21804:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21805:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21806:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21807:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21808:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd222;
        end
        21809:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd7;
        end
        21810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21812:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        21813:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        21814:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21815:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21816:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        21817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21818:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd124;
        end
        21819:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21820:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21821:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21822:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21823:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21824:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21825:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21826:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21827:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd139;
        end
        21828:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        21829:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        21830:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        21831:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21832:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21833:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21834:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21835:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21836:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21837:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21838:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        21839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21842:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        21843:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        21844:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21845:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21846:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21847:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21848:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21849:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21850:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21851:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        21852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21876:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd121;
        end
        21877:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21878:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21879:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21880:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21881:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21882:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21884:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd179;
        end
        21885:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd6;
        end
        21886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21890:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd56;
        end
        21891:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd232;
        end
        21892:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21893:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21894:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21895:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21896:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21897:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21898:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd224;
        end
        21899:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd39;
        end
        21900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21905:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd94;
        end
        21906:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21908:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21909:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21910:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21911:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21912:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21913:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21914:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21915:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21916:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21917:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd51;
        end
        21918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21924:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        21925:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21926:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21927:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21928:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21929:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21930:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21932:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        21933:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        21934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21946:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        21947:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21948:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21949:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21950:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21951:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21952:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21954:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        21955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21958:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd49;
        end
        21959:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        21960:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21961:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21962:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21963:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21964:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21965:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        21966:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd229;
        end
        21967:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd65;
        end
        21968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        21973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22020:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd22;
        end
        22021:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd232;
        end
        22022:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22023:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22024:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22025:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22026:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22027:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22028:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22029:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd80;
        end
        22030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22035:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        22036:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22037:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22038:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22039:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22040:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22041:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22042:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22043:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        22044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22045:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd7;
        end
        22046:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd185;
        end
        22047:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22048:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22049:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22050:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22051:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22052:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22053:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22054:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22055:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22056:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22057:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22058:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22059:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22060:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22061:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22062:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22063:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22064:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22065:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd19;
        end
        22066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22068:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        22069:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        22070:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22071:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22072:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        22073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22074:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd99;
        end
        22075:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22076:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22077:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22078:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22079:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22080:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22081:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22082:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22083:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd111;
        end
        22084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22085:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        22086:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        22087:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22088:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22089:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22090:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22091:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22092:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22093:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22094:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        22095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22098:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        22099:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        22100:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22101:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22102:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22103:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22104:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22105:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22106:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22107:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        22108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22132:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd92;
        end
        22133:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        22134:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22135:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22136:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22137:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22138:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22139:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22140:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd185;
        end
        22141:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd7;
        end
        22142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22146:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd63;
        end
        22147:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22148:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22149:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22150:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22151:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22152:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22153:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22154:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd210;
        end
        22155:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd26;
        end
        22156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22161:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd72;
        end
        22162:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd232;
        end
        22163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22164:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22165:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22166:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22167:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22168:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22169:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22170:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22171:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22172:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22173:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd27;
        end
        22174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22180:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        22181:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22182:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22183:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22185:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22186:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22188:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        22189:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        22190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22202:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        22203:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22204:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22205:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22206:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22207:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22208:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22210:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        22211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22214:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd42;
        end
        22215:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd227;
        end
        22216:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22217:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22218:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22219:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22220:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22221:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22222:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd230;
        end
        22223:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd70;
        end
        22224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22276:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd2;
        end
        22277:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd214;
        end
        22278:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22279:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22280:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22281:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22282:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22283:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22284:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22285:
        begin
            RED=8'd0;
            GRN=8'd90;
            BLU=8'd98;
        end
        22286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22291:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        22292:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22293:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22294:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22295:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22296:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22297:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22298:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22299:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        22300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22301:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd12;
        end
        22302:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd203;
        end
        22303:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22304:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22305:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22306:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22307:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22308:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22309:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22310:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22311:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22312:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22313:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22314:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22315:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22316:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22317:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22318:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22319:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22320:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22321:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd43;
        end
        22322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22324:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        22325:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        22326:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22327:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22328:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        22329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22330:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd69;
        end
        22331:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd231;
        end
        22332:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22333:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22334:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22335:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22336:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22337:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22338:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22339:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd85;
        end
        22340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22341:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        22342:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        22343:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22344:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22345:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22347:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22348:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22349:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22350:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        22351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22354:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        22355:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        22356:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22357:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22358:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22359:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22360:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22361:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22362:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22363:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        22364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22388:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd63;
        end
        22389:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        22390:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22391:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22393:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22394:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22396:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd190;
        end
        22397:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd8;
        end
        22398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22402:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd70;
        end
        22403:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22404:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22405:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22406:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22407:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22408:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22409:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22410:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd194;
        end
        22411:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd11;
        end
        22412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22417:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd46;
        end
        22418:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd232;
        end
        22419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22420:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22421:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22422:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22423:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22424:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22425:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22426:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22427:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22428:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd222;
        end
        22429:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd15;
        end
        22430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22436:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        22437:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22438:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22439:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22441:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22442:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22443:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22444:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        22445:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        22446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22458:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        22459:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22460:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22461:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22462:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22463:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22464:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22465:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22466:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        22467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd35;
        end
        22471:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd226;
        end
        22472:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22473:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22474:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22475:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22476:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22477:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22478:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        22479:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd75;
        end
        22480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22532:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd2;
        end
        22533:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd180;
        end
        22534:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22535:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22536:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22537:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22538:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22539:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22540:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22541:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd113;
        end
        22542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22547:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        22548:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22549:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22550:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22551:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22552:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22553:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22554:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22555:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        22556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22557:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd16;
        end
        22558:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd218;
        end
        22559:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22560:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22561:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd210;
        end
        22562:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd152;
        end
        22563:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd150;
        end
        22564:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd150;
        end
        22565:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd150;
        end
        22566:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd150;
        end
        22567:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd150;
        end
        22568:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd163;
        end
        22569:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd227;
        end
        22570:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22571:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22572:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22573:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22574:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22575:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22576:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22577:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd72;
        end
        22578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22580:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        22581:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        22582:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22583:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22584:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        22585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22586:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd42;
        end
        22587:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd231;
        end
        22588:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22589:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22590:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22591:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22592:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22593:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22594:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd229;
        end
        22595:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd66;
        end
        22596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22597:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        22598:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        22599:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22600:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22601:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22603:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22604:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22605:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22606:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        22607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22610:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        22611:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        22612:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22613:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22614:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22615:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22616:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22617:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22618:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22619:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        22620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22644:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd38;
        end
        22645:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd219;
        end
        22646:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22647:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22648:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22649:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22650:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22652:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd201;
        end
        22653:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd11;
        end
        22654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22658:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd84;
        end
        22659:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22660:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22661:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22662:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22663:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22664:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22665:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22666:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd168;
        end
        22667:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        22668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22673:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd30;
        end
        22674:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd225;
        end
        22675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22676:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22677:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22678:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22679:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22680:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22681:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22682:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22683:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22684:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd200;
        end
        22685:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd10;
        end
        22686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22692:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        22693:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22694:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22695:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22696:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22698:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22699:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22700:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        22701:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        22702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22714:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        22715:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22716:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22717:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22718:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22719:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22720:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22721:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22722:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        22723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd35;
        end
        22727:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd226;
        end
        22728:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22729:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22730:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22731:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22732:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22733:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22734:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22735:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd82;
        end
        22736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        22789:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd142;
        end
        22790:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22791:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22792:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22793:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22794:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22795:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22796:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22797:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd127;
        end
        22798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22803:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        22804:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22805:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22806:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22807:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22808:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22809:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22810:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22811:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        22812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22813:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd29;
        end
        22814:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd232;
        end
        22815:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22816:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22817:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd162;
        end
        22818:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd3;
        end
        22819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22824:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd33;
        end
        22825:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd217;
        end
        22826:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22827:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22828:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22829:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22830:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22831:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22832:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22833:
        begin
            RED=8'd0;
            GRN=8'd94;
            BLU=8'd100;
        end
        22834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22836:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        22837:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        22838:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22839:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22840:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        22841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd15;
        end
        22843:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd231;
        end
        22844:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22845:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22846:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22847:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22848:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22849:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22850:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd223;
        end
        22851:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd46;
        end
        22852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22853:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        22854:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        22855:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22856:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22857:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22859:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22860:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22861:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22862:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        22863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22866:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        22867:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        22868:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22869:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22870:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22871:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22872:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22873:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22874:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22875:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        22876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd16;
        end
        22901:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd202;
        end
        22902:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22903:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22904:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22905:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22906:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22908:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd213;
        end
        22909:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd13;
        end
        22910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22914:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd98;
        end
        22915:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22916:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22917:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22918:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22919:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22920:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22921:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22922:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd132;
        end
        22923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22929:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd21;
        end
        22930:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd209;
        end
        22931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22932:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22933:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22934:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22935:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22936:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22937:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22938:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22939:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22940:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd175;
        end
        22941:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd5;
        end
        22942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22948:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        22949:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22950:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22951:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22952:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22954:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22955:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22956:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        22957:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        22958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22970:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        22971:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22972:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22973:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22974:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22975:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22976:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22977:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22978:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        22979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd35;
        end
        22983:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd226;
        end
        22984:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22985:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22986:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22987:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22988:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22989:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22990:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        22991:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd88;
        end
        22992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        22997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23045:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd86;
        end
        23046:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        23047:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23048:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23049:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23050:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23051:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23052:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23053:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd143;
        end
        23054:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        23055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23059:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd205;
        end
        23060:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23061:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23062:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23063:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23064:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23065:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23066:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23067:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        23068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23069:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd64;
        end
        23070:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23071:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23072:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23073:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd133;
        end
        23074:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        23075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd21;
        end
        23081:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd211;
        end
        23082:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23083:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23084:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23085:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23086:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23087:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23088:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23089:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd129;
        end
        23090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23092:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        23093:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        23094:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23095:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23096:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        23097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23099:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd226;
        end
        23100:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23101:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23102:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23103:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23104:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23105:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23106:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd217;
        end
        23107:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd27;
        end
        23108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23109:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        23110:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        23111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23113:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23114:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23115:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23116:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23117:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23118:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        23119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23122:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        23123:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        23124:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23125:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23126:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23127:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23128:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23129:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23130:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23131:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        23132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23157:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd182;
        end
        23158:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23159:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23161:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23162:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23164:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd223;
        end
        23165:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd15;
        end
        23166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23170:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd110;
        end
        23171:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23172:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23173:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23174:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23175:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23176:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23177:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        23178:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd99;
        end
        23179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd13;
        end
        23186:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd193;
        end
        23187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23188:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23189:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23190:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23191:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23192:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23193:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23194:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23195:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23196:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd150;
        end
        23197:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        23198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23204:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        23205:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23206:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23207:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23208:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23210:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23211:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23212:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        23213:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        23214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23226:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        23227:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23228:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23229:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23230:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23231:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23232:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23233:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23234:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        23235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd35;
        end
        23239:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd226;
        end
        23240:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23241:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23242:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23243:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23244:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23245:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23246:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23247:
        begin
            RED=8'd0;
            GRN=8'd97;
            BLU=8'd106;
        end
        23248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23301:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd39;
        end
        23302:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd228;
        end
        23303:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23304:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23305:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23306:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23307:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23308:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23309:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd168;
        end
        23310:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd1;
        end
        23311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        23315:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd206;
        end
        23316:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23317:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23318:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23319:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23320:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23321:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23322:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23323:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        23324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23325:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd91;
        end
        23326:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23327:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23328:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23329:
        begin
            RED=8'd0;
            GRN=8'd95;
            BLU=8'd106;
        end
        23330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23337:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd198;
        end
        23338:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23339:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23340:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23341:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23342:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23343:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23344:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23345:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd146;
        end
        23346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23348:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        23349:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        23350:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23351:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23352:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        23353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23355:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd200;
        end
        23356:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23357:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23358:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23359:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23360:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23361:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23362:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd212;
        end
        23363:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd14;
        end
        23364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23365:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        23366:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        23367:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23368:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23369:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23370:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23371:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23372:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23373:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23374:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        23375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23378:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        23379:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        23380:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23381:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23382:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23383:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23384:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23385:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23386:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23387:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        23388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23413:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd141;
        end
        23414:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23415:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23417:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23418:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23420:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23421:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd22;
        end
        23422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23426:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd125;
        end
        23427:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23428:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23429:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23430:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23431:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23432:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23433:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        23434:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd55;
        end
        23435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd7;
        end
        23442:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd181;
        end
        23443:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23444:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23445:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23446:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23447:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23448:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23449:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23450:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23451:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23452:
        begin
            RED=8'd0;
            GRN=8'd116;
            BLU=8'd136;
        end
        23453:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        23454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23460:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        23461:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23462:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23463:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23464:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23465:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23466:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23467:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23468:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        23469:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        23470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23482:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        23483:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23484:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23485:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23486:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23487:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23488:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23489:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23490:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        23491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd35;
        end
        23495:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd226;
        end
        23496:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23497:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23498:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23499:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23500:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23501:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23502:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23503:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd120;
        end
        23504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd17;
        end
        23558:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd199;
        end
        23559:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23560:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23561:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23562:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23563:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23564:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23565:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd193;
        end
        23566:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd12;
        end
        23567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd16;
        end
        23571:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd211;
        end
        23572:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23573:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23574:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23575:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23576:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23577:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23578:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23579:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        23580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23581:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd115;
        end
        23582:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23583:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23584:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23585:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd77;
        end
        23586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23593:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd186;
        end
        23594:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23595:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23596:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23597:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23598:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23599:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23600:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23601:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd174;
        end
        23602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23604:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        23605:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        23606:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23607:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23608:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        23609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23611:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd172;
        end
        23612:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23613:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23614:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23615:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23616:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23617:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23618:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd195;
        end
        23619:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd0;
        end
        23620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23621:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        23622:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        23623:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23624:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23625:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23626:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23627:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23628:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23629:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23630:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        23631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23634:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        23635:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        23636:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23637:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23638:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23639:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23640:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23641:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23642:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23643:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        23644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23669:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd79;
        end
        23670:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        23671:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23673:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23674:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23676:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23677:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd57;
        end
        23678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23682:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd161;
        end
        23683:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23684:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23685:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23686:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23687:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23688:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23689:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd221;
        end
        23690:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd0;
        end
        23691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23698:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd157;
        end
        23699:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23700:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23701:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23702:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23703:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23704:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23705:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23706:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23707:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23708:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd109;
        end
        23709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23716:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        23717:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23718:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23719:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23720:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23721:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23722:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23723:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23724:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        23725:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        23726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23738:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        23739:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23740:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23741:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23742:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23743:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23744:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23745:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23746:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        23747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd35;
        end
        23751:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd226;
        end
        23752:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23753:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23754:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23755:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23756:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23757:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23758:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23759:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd120;
        end
        23760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23814:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd151;
        end
        23815:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23816:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23817:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23818:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23819:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23820:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23821:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd223;
        end
        23822:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd26;
        end
        23823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd28;
        end
        23827:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd216;
        end
        23828:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23829:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23830:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23831:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23832:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23833:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23834:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23835:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        23836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23837:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd137;
        end
        23838:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23839:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23840:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23841:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd56;
        end
        23842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23849:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd158;
        end
        23850:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23851:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23852:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23853:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23854:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23855:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23856:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23857:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd200;
        end
        23858:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd0;
        end
        23859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23860:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        23861:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        23862:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23863:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23864:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        23865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23867:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd134;
        end
        23868:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23869:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23870:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23871:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23872:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23873:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23874:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd167;
        end
        23875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23877:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        23878:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        23879:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23880:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23881:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23882:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23884:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23885:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23886:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        23887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23890:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        23891:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        23892:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23893:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23894:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23895:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23896:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23897:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23898:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23899:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        23900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd21;
        end
        23926:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd230;
        end
        23927:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23928:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23929:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23930:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23932:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23933:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd87;
        end
        23934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23938:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd190;
        end
        23939:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23940:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23941:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23942:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23943:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23944:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23945:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd180;
        end
        23946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23954:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd142;
        end
        23955:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23956:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23957:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23958:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23959:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23960:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23961:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23962:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23963:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23964:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd77;
        end
        23965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23972:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        23973:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23974:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23975:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23976:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23977:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23978:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23979:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23980:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        23981:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        23982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        23994:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        23995:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23996:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23997:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23998:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        23999:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24000:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24001:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24002:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        24003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd35;
        end
        24007:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd226;
        end
        24008:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24009:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24010:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24011:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24012:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24013:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24014:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24015:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd136;
        end
        24016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24070:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd74;
        end
        24071:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd230;
        end
        24072:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24073:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24074:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24075:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24076:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24077:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        24078:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd66;
        end
        24079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24082:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd49;
        end
        24083:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd223;
        end
        24084:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24085:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24086:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24087:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24088:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24089:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24090:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24091:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        24092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24093:
        begin
            RED=8'd0;
            GRN=8'd95;
            BLU=8'd167;
        end
        24094:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24095:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24096:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd222;
        end
        24097:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd41;
        end
        24098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24105:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd127;
        end
        24106:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24107:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24108:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24109:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24110:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24113:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd207;
        end
        24114:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd14;
        end
        24115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24116:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        24117:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        24118:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24119:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24120:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        24121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24123:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd122;
        end
        24124:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24125:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24126:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24127:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24128:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24129:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24130:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd152;
        end
        24131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24133:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        24134:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        24135:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24136:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24137:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24138:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24139:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24140:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24141:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24142:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        24143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24146:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        24147:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        24148:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24149:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24150:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24151:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24152:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24153:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24154:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24155:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        24156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        24182:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd189;
        end
        24183:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24185:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24186:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24188:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24189:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        24190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24194:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd216;
        end
        24195:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24196:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24197:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24198:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24199:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24200:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24201:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd102;
        end
        24202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24210:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd113;
        end
        24211:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24212:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24213:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24214:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24215:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24216:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24217:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24218:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24219:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd226;
        end
        24220:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd49;
        end
        24221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24228:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        24229:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24230:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24231:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24232:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24233:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24234:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24235:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24236:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        24237:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        24238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24250:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        24251:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24252:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24253:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24254:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24255:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24256:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24257:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24258:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        24259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd20;
        end
        24263:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        24264:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24265:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24266:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24267:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24268:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24269:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24270:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24271:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd150;
        end
        24272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24326:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd9;
        end
        24327:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd219;
        end
        24328:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24329:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24330:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24331:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24332:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24333:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24334:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd137;
        end
        24335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24338:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd100;
        end
        24339:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd231;
        end
        24340:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24341:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24342:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24343:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24344:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24345:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24347:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        24348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24349:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd194;
        end
        24350:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24351:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24352:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd210;
        end
        24353:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd25;
        end
        24354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24361:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd107;
        end
        24362:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24363:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24364:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24365:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24366:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24367:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24368:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24369:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd217;
        end
        24370:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd33;
        end
        24371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24372:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        24373:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        24374:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24375:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24376:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        24377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24379:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd96;
        end
        24380:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24381:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24382:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24383:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24384:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24385:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24386:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd118;
        end
        24387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24389:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        24390:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        24391:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24393:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24394:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24396:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24397:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24398:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        24399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24402:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        24403:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        24404:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24405:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24406:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24407:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24408:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24409:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24410:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24411:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        24412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24438:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd129;
        end
        24439:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24441:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24442:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24443:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24444:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24445:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd161;
        end
        24446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24449:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd40;
        end
        24450:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd225;
        end
        24451:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24452:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24453:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24454:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24455:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24456:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24457:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd38;
        end
        24458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24466:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd78;
        end
        24467:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        24468:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24469:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24470:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24471:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24472:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24473:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24474:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24475:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd221;
        end
        24476:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd41;
        end
        24477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24484:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        24485:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24486:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24487:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24488:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24489:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24490:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24491:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24492:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        24493:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        24494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24506:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        24507:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24508:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24509:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24510:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24511:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24512:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24513:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24514:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        24515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd19;
        end
        24519:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        24520:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24521:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24522:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24523:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24524:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24525:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24526:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24527:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd163;
        end
        24528:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd0;
        end
        24529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24583:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd158;
        end
        24584:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24585:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24586:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24587:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24588:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24589:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24590:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd209;
        end
        24591:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd27;
        end
        24592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24593:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd9;
        end
        24594:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd175;
        end
        24595:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24596:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24597:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24598:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24599:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24600:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24601:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24603:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        24604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd13;
        end
        24605:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd212;
        end
        24606:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24607:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24608:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd202;
        end
        24609:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd15;
        end
        24610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24617:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd82;
        end
        24618:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24619:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24620:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24621:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24622:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24623:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24624:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24625:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd226;
        end
        24626:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd52;
        end
        24627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24628:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        24629:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        24630:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24631:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24632:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        24633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24635:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd66;
        end
        24636:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        24637:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24638:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24639:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24640:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24641:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24642:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd91;
        end
        24643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24645:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        24646:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        24647:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24648:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24649:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24650:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24652:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24653:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24654:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        24655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24658:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        24659:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        24660:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24661:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24662:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24663:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24664:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24665:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24666:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24667:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd78;
        end
        24668:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24669:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24670:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24671:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24672:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24673:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24674:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24675:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24676:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24677:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24678:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd9;
        end
        24679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24694:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd50;
        end
        24695:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd226;
        end
        24696:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24698:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24699:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24700:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24701:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd208;
        end
        24702:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd24;
        end
        24703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24705:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd105;
        end
        24706:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd231;
        end
        24707:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24708:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24709:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24710:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24711:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24712:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd191;
        end
        24713:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd12;
        end
        24714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24722:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd65;
        end
        24723:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd229;
        end
        24724:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24725:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24726:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24727:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24728:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24729:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24730:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24731:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd211;
        end
        24732:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd26;
        end
        24733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24740:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        24741:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24742:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24743:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24744:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24745:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24746:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24747:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24748:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd218;
        end
        24749:
        begin
            RED=8'd0;
            GRN=8'd59;
            BLU=8'd66;
        end
        24750:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24751:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24752:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24753:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24754:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24755:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24756:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24757:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24758:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24759:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd41;
        end
        24760:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        24761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24762:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        24763:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24764:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24765:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24766:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24767:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24768:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24769:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24770:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        24771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        24775:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd223;
        end
        24776:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24777:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24778:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24779:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24780:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24781:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24782:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24783:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd175;
        end
        24784:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd0;
        end
        24785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24839:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd57;
        end
        24840:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd225;
        end
        24841:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24842:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24843:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24844:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24845:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24846:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd230;
        end
        24847:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd159;
        end
        24848:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd60;
        end
        24849:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd123;
        end
        24850:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd220;
        end
        24851:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24852:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24853:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24854:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24855:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24856:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24857:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24859:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        24860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd27;
        end
        24861:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd219;
        end
        24862:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24863:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24864:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd186;
        end
        24865:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd4;
        end
        24866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24873:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd55;
        end
        24874:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24875:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24876:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24877:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24878:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24879:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24880:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24881:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        24882:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd62;
        end
        24883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24884:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        24885:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        24886:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24887:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24888:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        24889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24891:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd41;
        end
        24892:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd226;
        end
        24893:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24894:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24895:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24896:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24897:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24898:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd74;
        end
        24899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24901:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        24902:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        24903:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24904:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24905:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24906:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24908:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24909:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24910:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        24911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24914:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        24915:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        24916:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24917:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24918:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24919:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24920:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24921:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24922:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24923:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd188;
        end
        24924:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24925:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24926:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24927:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24928:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24929:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24930:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24931:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24932:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24933:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        24934:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd39;
        end
        24935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24950:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd9;
        end
        24951:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd178;
        end
        24952:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24954:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24955:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24956:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24957:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd228;
        end
        24958:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd88;
        end
        24959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24960:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd12;
        end
        24961:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd176;
        end
        24962:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24963:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24964:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24965:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24966:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24967:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24968:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd117;
        end
        24969:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd2;
        end
        24970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24978:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd47;
        end
        24979:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd224;
        end
        24980:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24981:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24982:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24983:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24984:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24985:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24986:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24987:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd196;
        end
        24988:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd7;
        end
        24989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        24996:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        24997:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24998:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        24999:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25000:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25001:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25002:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25003:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25004:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd228;
        end
        25005:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd185;
        end
        25006:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25007:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25008:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25009:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25010:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25011:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25012:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25013:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25014:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25015:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd178;
        end
        25016:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd14;
        end
        25017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25018:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        25019:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25020:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25021:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25022:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25023:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25024:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25025:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25026:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        25027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25031:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        25032:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25033:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25034:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25035:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25036:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25037:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25038:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25039:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd193;
        end
        25040:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd12;
        end
        25041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25095:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd8;
        end
        25096:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd166;
        end
        25097:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25098:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25099:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25100:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25101:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25102:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25103:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd224;
        end
        25104:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd176;
        end
        25105:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd208;
        end
        25106:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25107:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25108:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25109:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25110:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25113:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25114:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25115:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        25116:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd45;
        end
        25117:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd224;
        end
        25118:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25119:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25120:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd161;
        end
        25121:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        25122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25129:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd35;
        end
        25130:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd232;
        end
        25131:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25132:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25133:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25134:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25135:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25136:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25137:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25138:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd89;
        end
        25139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25140:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        25141:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        25142:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25143:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25144:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        25145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25147:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd29;
        end
        25148:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd218;
        end
        25149:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25150:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25151:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25152:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25153:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25154:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd50;
        end
        25155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25157:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        25158:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        25159:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25161:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25162:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25164:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25165:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25166:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        25167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25170:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        25171:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        25172:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25173:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25174:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25175:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25176:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25177:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25178:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25179:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25180:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25181:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25182:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25183:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25185:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25186:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25188:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25189:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25190:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd51;
        end
        25191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25207:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd94;
        end
        25208:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd228;
        end
        25209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25210:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25211:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25212:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25213:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25214:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd182;
        end
        25215:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd67;
        end
        25216:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd117;
        end
        25217:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd220;
        end
        25218:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25219:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25220:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25221:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25222:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25223:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd206;
        end
        25224:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd34;
        end
        25225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25234:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd34;
        end
        25235:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd220;
        end
        25236:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25237:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25238:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25239:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25240:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25241:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25242:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25243:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd174;
        end
        25244:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd0;
        end
        25245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25252:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        25253:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25254:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25255:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25256:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25257:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25258:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25259:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25260:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25261:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25262:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25263:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25264:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25265:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25266:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25267:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25268:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25269:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25270:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25271:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25272:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd19;
        end
        25273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25274:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        25275:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25276:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25277:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25278:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25279:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25280:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25281:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25282:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        25283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25287:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd200;
        end
        25288:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25289:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25290:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25291:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25292:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25293:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25294:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25295:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd205;
        end
        25296:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd21;
        end
        25297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25352:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd74;
        end
        25353:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd221;
        end
        25354:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25355:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25356:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25357:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25358:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25359:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25360:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25361:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25362:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25363:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25364:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25365:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25366:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd229;
        end
        25367:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd227;
        end
        25368:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25369:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25370:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25371:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        25372:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd66;
        end
        25373:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd229;
        end
        25374:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25375:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25376:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd132;
        end
        25377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25385:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd16;
        end
        25386:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd225;
        end
        25387:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25388:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25389:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25390:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25391:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25393:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25394:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd120;
        end
        25395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25396:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        25397:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        25398:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25399:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25400:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        25401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25403:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd20;
        end
        25404:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd205;
        end
        25405:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25406:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25407:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25408:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25409:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd226;
        end
        25410:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd25;
        end
        25411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25413:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        25414:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        25415:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25417:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25418:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25420:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25421:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25422:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        25423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25426:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        25427:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        25428:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25429:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25430:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25431:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25432:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25433:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25434:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25435:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25436:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25437:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25438:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25439:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25441:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25442:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25443:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25444:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25445:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25446:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd51;
        end
        25447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25463:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd25;
        end
        25464:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd187;
        end
        25465:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25466:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25467:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25468:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25469:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25470:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        25471:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd175;
        end
        25472:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd207;
        end
        25473:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25474:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25475:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25476:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25477:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25478:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25479:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd123;
        end
        25480:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        25481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd13;
        end
        25491:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd213;
        end
        25492:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25493:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25494:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25495:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25496:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25497:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25498:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25499:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd156;
        end
        25500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25508:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        25509:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25510:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25511:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25512:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25513:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25514:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25515:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25516:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25517:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25518:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25519:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25520:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25521:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25522:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25523:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25524:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25525:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25526:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25527:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25528:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd19;
        end
        25529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25530:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        25531:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25532:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25533:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25534:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25535:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25536:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25537:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25538:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        25539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25543:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd187;
        end
        25544:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25545:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25546:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25547:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25548:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25549:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25550:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25551:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd217;
        end
        25552:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd31;
        end
        25553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25608:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd14;
        end
        25609:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd149;
        end
        25610:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        25611:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25612:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25613:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25614:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25615:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25616:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25617:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25618:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25619:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25620:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25621:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25622:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd181;
        end
        25623:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd198;
        end
        25624:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25625:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25626:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25627:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        25628:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd94;
        end
        25629:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        25630:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25631:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25632:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd107;
        end
        25633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25641:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd5;
        end
        25642:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd214;
        end
        25643:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25644:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25645:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25646:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25647:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25648:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25649:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25650:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd140;
        end
        25651:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd0;
        end
        25652:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        25653:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        25654:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25655:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25656:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        25657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd8;
        end
        25660:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd186;
        end
        25661:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25662:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25663:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25664:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25665:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd215;
        end
        25666:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd13;
        end
        25667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25669:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        25670:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        25671:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25673:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25674:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25676:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25677:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25678:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        25679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25682:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        25683:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        25684:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25685:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25686:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25687:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25688:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25689:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25690:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25691:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25692:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25693:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25694:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25695:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25696:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25698:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25699:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25700:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25701:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25702:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd51;
        end
        25703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25720:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd99;
        end
        25721:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd222;
        end
        25722:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25723:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25724:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25725:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25726:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25727:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25728:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25729:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25730:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25731:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25732:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25733:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25734:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd196;
        end
        25735:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd36;
        end
        25736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25747:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd196;
        end
        25748:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25749:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25750:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25751:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25752:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25753:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25754:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25755:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd134;
        end
        25756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25764:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        25765:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25766:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25767:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25768:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25769:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25770:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25771:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25772:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25773:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25774:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25775:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25776:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25777:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25778:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25779:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25780:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25781:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25782:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25783:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25784:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd19;
        end
        25785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25786:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        25787:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25788:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25789:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25790:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25791:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25792:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25793:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25794:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        25795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25799:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd173;
        end
        25800:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25801:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25802:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25803:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25804:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25805:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25806:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25807:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        25808:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd57;
        end
        25809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25865:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd47;
        end
        25866:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd182;
        end
        25867:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        25868:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25869:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25870:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25871:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25872:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25873:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25874:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25875:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25876:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25877:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd206;
        end
        25878:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd80;
        end
        25879:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd153;
        end
        25880:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25881:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25882:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25883:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        25884:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd126;
        end
        25885:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25886:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25887:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25888:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd85;
        end
        25889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25897:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd4;
        end
        25898:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd196;
        end
        25899:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25900:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25901:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25902:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25903:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25904:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25905:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25906:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd159;
        end
        25907:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd2;
        end
        25908:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        25909:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        25910:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25911:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25912:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        25913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25916:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd168;
        end
        25917:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25918:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25919:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25920:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25921:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd199;
        end
        25922:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd10;
        end
        25923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25925:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        25926:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        25927:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25928:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25929:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25930:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25932:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25933:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25934:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        25935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25938:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        25939:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        25940:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25941:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25942:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25943:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25944:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25945:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25946:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25947:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25948:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25949:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25950:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25951:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25952:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25954:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25955:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25956:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25957:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25958:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd51;
        end
        25959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25976:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd22;
        end
        25977:
        begin
            RED=8'd0;
            GRN=8'd94;
            BLU=8'd154;
        end
        25978:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        25979:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25980:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25981:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25982:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25983:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25984:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25985:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25986:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25987:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25988:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        25989:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd213;
        end
        25990:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd99;
        end
        25991:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd2;
        end
        25992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        25999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26003:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd176;
        end
        26004:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26005:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26006:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26007:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26008:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26009:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26010:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26011:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd104;
        end
        26012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26020:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        26021:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26022:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26023:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26024:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26025:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26026:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26027:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26028:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26029:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26030:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26031:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26032:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26033:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26034:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26035:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26036:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26037:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26038:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26039:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26040:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd19;
        end
        26041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26042:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        26043:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26044:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26045:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26046:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26047:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26048:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26049:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26050:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        26051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26055:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd150;
        end
        26056:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26057:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26058:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26059:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26060:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26061:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26062:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26063:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26064:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd92;
        end
        26065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26122:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd70;
        end
        26123:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd187;
        end
        26124:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd231;
        end
        26125:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26126:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26127:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26128:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26129:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26130:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26131:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26132:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd212;
        end
        26133:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd118;
        end
        26134:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        26135:
        begin
            RED=8'd0;
            GRN=8'd59;
            BLU=8'd117;
        end
        26136:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        26137:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26138:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26139:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd2;
        end
        26140:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd149;
        end
        26141:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26142:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26143:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26144:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd59;
        end
        26145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        26154:
        begin
            RED=8'd0;
            GRN=8'd94;
            BLU=8'd168;
        end
        26155:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26156:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26157:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26158:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26159:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26161:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26162:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd184;
        end
        26163:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd8;
        end
        26164:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd74;
        end
        26165:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        26166:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26167:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26168:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd23;
        end
        26169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26172:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd151;
        end
        26173:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26174:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26175:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26176:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26177:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd174;
        end
        26178:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd5;
        end
        26179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26181:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd38;
        end
        26182:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        26183:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26185:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26186:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26187:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26188:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26189:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26190:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd28;
        end
        26191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26194:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd62;
        end
        26195:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd229;
        end
        26196:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26197:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26198:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26199:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26200:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26201:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26202:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26203:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26204:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26205:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26206:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26207:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26208:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26210:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26211:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26212:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26213:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26214:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd51;
        end
        26215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26233:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd44;
        end
        26234:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd167;
        end
        26235:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd228;
        end
        26236:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26237:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26238:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26239:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26240:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26241:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26242:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26243:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26244:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd214;
        end
        26245:
        begin
            RED=8'd0;
            GRN=8'd97;
            BLU=8'd129;
        end
        26246:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd8;
        end
        26247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26259:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd157;
        end
        26260:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26261:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26262:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26263:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26264:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26265:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26266:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26267:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd73;
        end
        26268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26276:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd91;
        end
        26277:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26278:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26279:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26280:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26281:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26282:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26283:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26284:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26285:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26286:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26287:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26288:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26289:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26290:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26291:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26292:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26293:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26294:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26295:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26296:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd19;
        end
        26297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26298:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd182;
        end
        26299:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26300:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26301:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26302:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26303:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26304:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26305:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26306:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd163;
        end
        26307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26311:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        26312:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26313:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26314:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26315:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26316:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26317:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26318:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26319:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26320:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd130;
        end
        26321:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        26322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26379:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd64;
        end
        26380:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd182;
        end
        26381:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd210;
        end
        26382:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd224;
        end
        26383:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26384:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26385:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26386:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd225;
        end
        26387:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd199;
        end
        26388:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd129;
        end
        26389:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd8;
        end
        26390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26391:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd74;
        end
        26392:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd182;
        end
        26393:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26394:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26395:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd2;
        end
        26396:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd125;
        end
        26397:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26398:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26399:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd181;
        end
        26400:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd30;
        end
        26401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26410:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd112;
        end
        26411:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26412:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26413:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26414:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26415:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26416:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26417:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26418:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd158;
        end
        26419:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd11;
        end
        26420:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd58;
        end
        26421:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd182;
        end
        26422:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26423:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26424:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd18;
        end
        26425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26428:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd103;
        end
        26429:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26430:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26431:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26432:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26433:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd119;
        end
        26434:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd0;
        end
        26435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26437:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd30;
        end
        26438:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd176;
        end
        26439:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26440:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26441:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26442:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26443:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26444:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26445:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26446:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd22;
        end
        26447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26450:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd49;
        end
        26451:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd179;
        end
        26452:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26453:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26454:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26455:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26456:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26457:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26458:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26459:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26460:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26461:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26462:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26463:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26464:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26465:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26466:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26467:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26468:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26469:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26470:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd40;
        end
        26471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26490:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd31;
        end
        26491:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd173;
        end
        26492:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd205;
        end
        26493:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd225;
        end
        26494:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        26495:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26496:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        26497:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd230;
        end
        26498:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd219;
        end
        26499:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd193;
        end
        26500:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd133;
        end
        26501:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd0;
        end
        26502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26515:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd105;
        end
        26516:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26517:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26518:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26519:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26520:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26521:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26522:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd181;
        end
        26523:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd42;
        end
        26524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26532:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd71;
        end
        26533:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26534:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26535:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26536:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26537:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26538:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26539:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26540:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26541:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26542:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26543:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26544:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26545:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26546:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26547:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26548:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26549:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26550:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26551:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26552:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd15;
        end
        26553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26554:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd143;
        end
        26555:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26556:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26557:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26558:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26559:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26560:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26561:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26562:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd128;
        end
        26563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26567:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd78;
        end
        26568:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26569:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26570:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26571:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26572:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26573:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26574:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26575:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        26576:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd138;
        end
        26577:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd1;
        end
        26578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26636:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd10;
        end
        26637:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd112;
        end
        26638:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd170;
        end
        26639:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd201;
        end
        26640:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd201;
        end
        26641:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd201;
        end
        26642:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd172;
        end
        26643:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd68;
        end
        26644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd8;
        end
        26748:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd93;
        end
        26749:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd173;
        end
        26750:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd201;
        end
        26751:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd201;
        end
        26752:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd201;
        end
        26753:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd191;
        end
        26754:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd150;
        end
        26755:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd43;
        end
        26756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        26999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        27999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        28999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        29999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        30999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31281:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd24;
        end
        31282:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd30;
        end
        31283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31294:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd29;
        end
        31295:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd25;
        end
        31296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31358:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd12;
        end
        31359:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd43;
        end
        31360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31530:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd14;
        end
        31531:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd143;
        end
        31532:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd176;
        end
        31533:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd161;
        end
        31534:
        begin
            RED=8'd0;
            GRN=8'd33;
            BLU=8'd32;
        end
        31535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31536:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd140;
        end
        31537:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd183;
        end
        31538:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd121;
        end
        31539:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd39;
        end
        31540:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd176;
        end
        31541:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd134;
        end
        31542:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd2;
        end
        31543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31549:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd161;
        end
        31550:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd184;
        end
        31551:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd98;
        end
        31552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31559:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd156;
        end
        31560:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd176;
        end
        31561:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd176;
        end
        31562:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd176;
        end
        31563:
        begin
            RED=8'd0;
            GRN=8'd116;
            BLU=8'd167;
        end
        31564:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd36;
        end
        31565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd14;
        end
        31586:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd19;
        end
        31587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31593:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd18;
        end
        31594:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd15;
        end
        31595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31606:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd91;
        end
        31607:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd176;
        end
        31608:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd176;
        end
        31609:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd176;
        end
        31610:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd176;
        end
        31611:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd104;
        end
        31612:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd0;
        end
        31613:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd89;
        end
        31614:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd179;
        end
        31615:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd175;
        end
        31616:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd0;
        end
        31617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31633:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd55;
        end
        31634:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd176;
        end
        31635:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd170;
        end
        31636:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd34;
        end
        31637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31651:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd79;
        end
        31652:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd176;
        end
        31653:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd96;
        end
        31654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        31786:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd107;
        end
        31787:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd218;
        end
        31788:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd157;
        end
        31789:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd181;
        end
        31790:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd124;
        end
        31791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31792:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        31793:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31794:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        31795:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd82;
        end
        31796:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd232;
        end
        31797:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd196;
        end
        31798:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd3;
        end
        31799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31805:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        31806:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31807:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd120;
        end
        31808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31815:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        31816:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31817:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31818:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31819:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd228;
        end
        31820:
        begin
            RED=8'd0;
            GRN=8'd122;
            BLU=8'd156;
        end
        31821:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd10;
        end
        31822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd6;
        end
        31841:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd125;
        end
        31842:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd84;
        end
        31843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd10;
        end
        31849:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd140;
        end
        31850:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd65;
        end
        31851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31862:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        31863:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31864:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31865:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31866:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31867:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd201;
        end
        31868:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd53;
        end
        31869:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        31870:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31871:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        31872:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd0;
        end
        31873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31889:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd93;
        end
        31890:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        31891:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd228;
        end
        31892:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd61;
        end
        31893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31898:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd113;
        end
        31899:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd145;
        end
        31900:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd21;
        end
        31901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31907:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd134;
        end
        31908:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        31909:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd148;
        end
        31910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        31957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32041:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd18;
        end
        32042:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd198;
        end
        32043:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32044:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd56;
        end
        32045:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd108;
        end
        32046:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd198;
        end
        32047:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd0;
        end
        32048:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        32049:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32050:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        32051:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd70;
        end
        32052:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        32053:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd189;
        end
        32054:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd2;
        end
        32055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32061:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        32062:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32063:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd120;
        end
        32064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32071:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        32072:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32073:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd202;
        end
        32074:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd154;
        end
        32075:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32076:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd222;
        end
        32077:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd59;
        end
        32078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32093:
        begin
            RED=8'd38;
            GRN=8'd54;
            BLU=8'd58;
        end
        32094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        32096:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd117;
        end
        32097:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd209;
        end
        32098:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        32099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32103:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd9;
        end
        32104:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd126;
        end
        32105:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd217;
        end
        32106:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        32107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32118:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        32119:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32120:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd227;
        end
        32121:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd139;
        end
        32122:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd222;
        end
        32123:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32124:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd122;
        end
        32125:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd118;
        end
        32126:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32127:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        32128:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd0;
        end
        32129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32145:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd119;
        end
        32146:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32147:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        32148:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd88;
        end
        32149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32153:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd20;
        end
        32154:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd195;
        end
        32155:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        32156:
        begin
            RED=8'd0;
            GRN=8'd59;
            BLU=8'd58;
        end
        32157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32163:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd122;
        end
        32164:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        32165:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd140;
        end
        32166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32297:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd67;
        end
        32298:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        32299:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd220;
        end
        32300:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd9;
        end
        32301:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd58;
        end
        32302:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd220;
        end
        32303:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd25;
        end
        32304:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        32305:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32306:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        32307:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd25;
        end
        32308:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd113;
        end
        32309:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd86;
        end
        32310:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        32311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32317:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        32318:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32319:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd120;
        end
        32320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32327:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        32328:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32329:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        32330:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd66;
        end
        32331:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd225;
        end
        32332:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32333:
        begin
            RED=8'd0;
            GRN=8'd95;
            BLU=8'd105;
        end
        32334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32349:
        begin
            RED=8'd31;
            GRN=8'd44;
            BLU=8'd47;
        end
        32350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32351:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd2;
        end
        32352:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd205;
        end
        32353:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32354:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        32355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32359:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd19;
        end
        32360:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd212;
        end
        32361:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32362:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        32363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32374:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        32375:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32376:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        32377:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd59;
        end
        32378:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd197;
        end
        32379:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32380:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd169;
        end
        32381:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd121;
        end
        32382:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32383:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        32384:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd0;
        end
        32385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32401:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd142;
        end
        32402:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32403:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32404:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd111;
        end
        32405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32409:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd38;
        end
        32410:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd218;
        end
        32411:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32412:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd77;
        end
        32413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32419:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd51;
        end
        32420:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd113;
        end
        32421:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd62;
        end
        32422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32553:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd127;
        end
        32554:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32555:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd196;
        end
        32556:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd6;
        end
        32557:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd43;
        end
        32558:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd218;
        end
        32559:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd54;
        end
        32560:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        32561:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32562:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        32563:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd0;
        end
        32564:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd5;
        end
        32565:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd29;
        end
        32566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        32567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32573:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        32574:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32575:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd120;
        end
        32576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32583:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        32584:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32585:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        32586:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd31;
        end
        32587:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd214;
        end
        32588:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32589:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd127;
        end
        32590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32607:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd2;
        end
        32608:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        32609:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32610:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        32611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32615:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        32616:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        32617:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32618:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        32619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32630:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        32631:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32632:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        32633:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        32634:
        begin
            RED=8'd0;
            GRN=8'd95;
            BLU=8'd167;
        end
        32635:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32636:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd196;
        end
        32637:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd127;
        end
        32638:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32639:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        32640:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd0;
        end
        32641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32657:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd166;
        end
        32658:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32659:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32660:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd132;
        end
        32661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32665:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd42;
        end
        32666:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd215;
        end
        32667:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd224;
        end
        32668:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd64;
        end
        32669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32676:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd10;
        end
        32677:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd26;
        end
        32678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32680:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd16;
        end
        32681:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd19;
        end
        32682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32809:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd173;
        end
        32810:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32811:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd176;
        end
        32812:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd3;
        end
        32813:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd38;
        end
        32814:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd216;
        end
        32815:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd57;
        end
        32816:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        32817:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32818:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        32819:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd39;
        end
        32820:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd89;
        end
        32821:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd121;
        end
        32822:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd3;
        end
        32823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32824:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd24;
        end
        32825:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd78;
        end
        32826:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd82;
        end
        32827:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd43;
        end
        32828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32829:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        32830:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32831:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd120;
        end
        32832:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd8;
        end
        32833:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd73;
        end
        32834:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd25;
        end
        32835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32839:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        32840:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32841:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        32842:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd27;
        end
        32843:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd210;
        end
        32844:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32845:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd131;
        end
        32846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32847:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd20;
        end
        32848:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd77;
        end
        32849:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd80;
        end
        32850:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd38;
        end
        32851:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        32852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32853:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd47;
        end
        32854:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd82;
        end
        32855:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd78;
        end
        32856:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd20;
        end
        32857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32859:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd45;
        end
        32860:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd82;
        end
        32861:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd74;
        end
        32862:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd15;
        end
        32863:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd50;
        end
        32864:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd224;
        end
        32865:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32866:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd154;
        end
        32867:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd33;
        end
        32868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32871:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd72;
        end
        32872:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd225;
        end
        32873:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32874:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd138;
        end
        32875:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd25;
        end
        32876:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd4;
        end
        32877:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd63;
        end
        32878:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd82;
        end
        32879:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd79;
        end
        32880:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd27;
        end
        32881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32886:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        32887:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32888:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        32889:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        32890:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd151;
        end
        32891:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32892:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd210;
        end
        32893:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd131;
        end
        32894:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32895:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        32896:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd0;
        end
        32897:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd28;
        end
        32898:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd76;
        end
        32899:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd82;
        end
        32900:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd76;
        end
        32901:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd25;
        end
        32902:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd49;
        end
        32903:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd82;
        end
        32904:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd78;
        end
        32905:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd9;
        end
        32906:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd15;
        end
        32907:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd79;
        end
        32908:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd3;
        end
        32909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32913:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd195;
        end
        32914:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32915:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        32916:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd159;
        end
        32917:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd0;
        end
        32918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32919:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd15;
        end
        32920:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd74;
        end
        32921:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd109;
        end
        32922:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd216;
        end
        32923:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd157;
        end
        32924:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd31;
        end
        32925:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd13;
        end
        32926:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd70;
        end
        32927:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd82;
        end
        32928:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd79;
        end
        32929:
        begin
            RED=8'd0;
            GRN=8'd33;
            BLU=8'd41;
        end
        32930:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        32931:
        begin
            RED=8'd0;
            GRN=8'd33;
            BLU=8'd57;
        end
        32932:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd96;
        end
        32933:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd99;
        end
        32934:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        32935:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd78;
        end
        32936:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd105;
        end
        32937:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd85;
        end
        32938:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd77;
        end
        32939:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd82;
        end
        32940:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd16;
        end
        32941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        32981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd7;
        end
        33065:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd203;
        end
        33066:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33067:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd160;
        end
        33068:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd1;
        end
        33069:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd32;
        end
        33070:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd175;
        end
        33071:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd35;
        end
        33072:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        33073:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33074:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        33075:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        33076:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33077:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        33078:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd4;
        end
        33079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd8;
        end
        33080:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd109;
        end
        33081:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd219;
        end
        33082:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd199;
        end
        33083:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd148;
        end
        33084:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd9;
        end
        33085:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        33086:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33087:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd120;
        end
        33088:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd38;
        end
        33089:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd208;
        end
        33090:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd54;
        end
        33091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33095:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        33096:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33097:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        33098:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd29;
        end
        33099:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd212;
        end
        33100:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33101:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd112;
        end
        33102:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        33103:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd91;
        end
        33104:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd223;
        end
        33105:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd218;
        end
        33106:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd140;
        end
        33107:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd6;
        end
        33108:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd20;
        end
        33109:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd161;
        end
        33110:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd195;
        end
        33111:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd208;
        end
        33112:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd92;
        end
        33113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33114:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd10;
        end
        33115:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd157;
        end
        33116:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd223;
        end
        33117:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd214;
        end
        33118:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd74;
        end
        33119:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd101;
        end
        33120:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd228;
        end
        33121:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33122:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd199;
        end
        33123:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd69;
        end
        33124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33127:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd124;
        end
        33128:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd229;
        end
        33129:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33130:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd193;
        end
        33131:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd51;
        end
        33132:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd39;
        end
        33133:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd193;
        end
        33134:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd216;
        end
        33135:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd227;
        end
        33136:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd116;
        end
        33137:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd1;
        end
        33138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33142:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        33143:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33144:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        33145:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        33146:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd151;
        end
        33147:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33148:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd210;
        end
        33149:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd131;
        end
        33150:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33151:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        33152:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd5;
        end
        33153:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd112;
        end
        33154:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd189;
        end
        33155:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd209;
        end
        33156:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd220;
        end
        33157:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd106;
        end
        33158:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd127;
        end
        33159:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        33160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd225;
        end
        33161:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd32;
        end
        33162:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd50;
        end
        33163:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd216;
        end
        33164:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd7;
        end
        33165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd5;
        end
        33169:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd218;
        end
        33170:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33171:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33172:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd180;
        end
        33173:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd2;
        end
        33174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        33175:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd82;
        end
        33176:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd215;
        end
        33177:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd225;
        end
        33178:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        33179:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd87;
        end
        33180:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd0;
        end
        33181:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd70;
        end
        33182:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd191;
        end
        33183:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd195;
        end
        33184:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd228;
        end
        33185:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd149;
        end
        33186:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd11;
        end
        33187:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        33188:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33189:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        33190:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        33191:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        33192:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33193:
        begin
            RED=8'd0;
            GRN=8'd139;
            BLU=8'd179;
        end
        33194:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd223;
        end
        33195:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33196:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd72;
        end
        33197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33320:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd28;
        end
        33321:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd214;
        end
        33322:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33323:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd146;
        end
        33324:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        33325:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd12;
        end
        33326:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd54;
        end
        33327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33328:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        33329:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33330:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        33331:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        33332:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33333:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        33334:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd4;
        end
        33335:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd46;
        end
        33336:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd221;
        end
        33337:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd208;
        end
        33338:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd97;
        end
        33339:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd217;
        end
        33340:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd36;
        end
        33341:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        33342:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33343:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd120;
        end
        33344:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd95;
        end
        33345:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd196;
        end
        33346:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd10;
        end
        33347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33351:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        33352:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33353:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        33354:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd47;
        end
        33355:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd221;
        end
        33356:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd228;
        end
        33357:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd77;
        end
        33358:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd13;
        end
        33359:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd191;
        end
        33360:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd227;
        end
        33361:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd179;
        end
        33362:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd224;
        end
        33363:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd35;
        end
        33364:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd89;
        end
        33365:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd232;
        end
        33366:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd88;
        end
        33367:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd157;
        end
        33368:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd193;
        end
        33369:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd3;
        end
        33370:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd56;
        end
        33371:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33372:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd184;
        end
        33373:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd222;
        end
        33374:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd169;
        end
        33375:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd7;
        end
        33376:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        33377:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33378:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        33379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33383:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        33384:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        33385:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33386:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        33387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33388:
        begin
            RED=8'd0;
            GRN=8'd69;
            BLU=8'd129;
        end
        33389:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33390:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd164;
        end
        33391:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd230;
        end
        33392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd222;
        end
        33393:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd18;
        end
        33394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33398:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        33399:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33400:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        33401:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        33402:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd156;
        end
        33403:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33404:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd205;
        end
        33405:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd130;
        end
        33406:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33407:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        33408:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd21;
        end
        33409:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd205;
        end
        33410:
        begin
            RED=8'd0;
            GRN=8'd95;
            BLU=8'd107;
        end
        33411:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd138;
        end
        33412:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33413:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd197;
        end
        33414:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd93;
        end
        33415:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd231;
        end
        33416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33417:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd57;
        end
        33418:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd80;
        end
        33419:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd187;
        end
        33420:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd4;
        end
        33421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd23;
        end
        33425:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd225;
        end
        33426:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd221;
        end
        33427:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33428:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd193;
        end
        33429:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd12;
        end
        33430:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd13;
        end
        33431:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd195;
        end
        33432:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd228;
        end
        33433:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd192;
        end
        33434:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        33435:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd186;
        end
        33436:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd8;
        end
        33437:
        begin
            RED=8'd0;
            GRN=8'd90;
            BLU=8'd166;
        end
        33438:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd160;
        end
        33439:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd85;
        end
        33440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33441:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33442:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd38;
        end
        33443:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        33444:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33445:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        33446:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        33447:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        33448:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33449:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd228;
        end
        33450:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd225;
        end
        33451:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33452:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd145;
        end
        33453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33576:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd36;
        end
        33577:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd218;
        end
        33578:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33579:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd146;
        end
        33580:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        33581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33584:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        33585:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33586:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        33587:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        33588:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33589:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        33590:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd4;
        end
        33591:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd118;
        end
        33592:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33593:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd173;
        end
        33594:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd36;
        end
        33595:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd226;
        end
        33596:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd51;
        end
        33597:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        33598:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33599:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd121;
        end
        33600:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd167;
        end
        33601:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd132;
        end
        33602:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        33603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33607:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        33608:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33609:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd187;
        end
        33610:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd115;
        end
        33611:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33612:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd198;
        end
        33613:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd24;
        end
        33614:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd55;
        end
        33615:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33616:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd205;
        end
        33617:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd132;
        end
        33618:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33619:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd100;
        end
        33620:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd153;
        end
        33621:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33622:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd68;
        end
        33623:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd91;
        end
        33624:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd210;
        end
        33625:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd18;
        end
        33626:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd140;
        end
        33627:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33628:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd125;
        end
        33629:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd212;
        end
        33630:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd217;
        end
        33631:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd31;
        end
        33632:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        33633:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33634:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        33635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33639:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        33640:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        33641:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33642:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        33643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        33644:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd199;
        end
        33645:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33646:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd119;
        end
        33647:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd217;
        end
        33648:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33649:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd80;
        end
        33650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33654:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        33655:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33656:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        33657:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd48;
        end
        33658:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd184;
        end
        33659:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33660:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd180;
        end
        33661:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd124;
        end
        33662:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33663:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        33664:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd37;
        end
        33665:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        33666:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd53;
        end
        33667:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd104;
        end
        33668:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33669:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd205;
        end
        33670:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd79;
        end
        33671:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd229;
        end
        33672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33673:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd86;
        end
        33674:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd121;
        end
        33675:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd158;
        end
        33676:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd2;
        end
        33677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33680:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd40;
        end
        33681:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd213;
        end
        33682:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd173;
        end
        33683:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33684:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd210;
        end
        33685:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd24;
        end
        33686:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd41;
        end
        33687:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd232;
        end
        33688:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd222;
        end
        33689:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd119;
        end
        33690:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        33691:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd221;
        end
        33692:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd42;
        end
        33693:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd202;
        end
        33694:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd113;
        end
        33695:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd45;
        end
        33696:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33698:
        begin
            RED=8'd0;
            GRN=8'd59;
            BLU=8'd54;
        end
        33699:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        33700:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33701:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        33702:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        33703:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        33704:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33705:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd209;
        end
        33706:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd193;
        end
        33707:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33708:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        33709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33832:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd36;
        end
        33833:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd218;
        end
        33834:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33835:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd146;
        end
        33836:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        33837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33840:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        33841:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33842:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        33843:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        33844:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33845:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        33846:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd4;
        end
        33847:
        begin
            RED=8'd0;
            GRN=8'd90;
            BLU=8'd158;
        end
        33848:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33849:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd148;
        end
        33850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd21;
        end
        33851:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd228;
        end
        33852:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd57;
        end
        33853:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        33854:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33855:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd125;
        end
        33856:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd232;
        end
        33857:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd78;
        end
        33858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33863:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        33864:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33865:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd231;
        end
        33866:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd230;
        end
        33867:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33868:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd66;
        end
        33869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33870:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd95;
        end
        33871:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33872:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd193;
        end
        33873:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd119;
        end
        33874:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33875:
        begin
            RED=8'd0;
            GRN=8'd122;
            BLU=8'd149;
        end
        33876:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd183;
        end
        33877:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33878:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd156;
        end
        33879:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd56;
        end
        33880:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd138;
        end
        33881:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd18;
        end
        33882:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd180;
        end
        33883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33884:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd112;
        end
        33885:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd199;
        end
        33886:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33887:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd60;
        end
        33888:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        33889:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33890:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        33891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33895:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        33896:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        33897:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33898:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        33899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd20;
        end
        33900:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd225;
        end
        33901:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33902:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd102;
        end
        33903:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd195;
        end
        33904:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33905:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd125;
        end
        33906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33910:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        33911:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33912:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        33913:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd89;
        end
        33914:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd221;
        end
        33915:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33916:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd137;
        end
        33917:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd118;
        end
        33918:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33919:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        33920:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd36;
        end
        33921:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd219;
        end
        33922:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd53;
        end
        33923:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd120;
        end
        33924:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33925:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd212;
        end
        33926:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd61;
        end
        33927:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd224;
        end
        33928:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33929:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd113;
        end
        33930:
        begin
            RED=8'd0;
            GRN=8'd82;
            BLU=8'd147;
        end
        33931:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd115;
        end
        33932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33936:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd66;
        end
        33937:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd210;
        end
        33938:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd136;
        end
        33939:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33940:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd224;
        end
        33941:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd35;
        end
        33942:
        begin
            RED=8'd0;
            GRN=8'd26;
            BLU=8'd76;
        end
        33943:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33944:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd220;
        end
        33945:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd89;
        end
        33946:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd232;
        end
        33947:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33948:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd56;
        end
        33949:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd197;
        end
        33950:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd111;
        end
        33951:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd62;
        end
        33952:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33954:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd68;
        end
        33955:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        33956:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33957:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        33958:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        33959:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        33960:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33961:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd167;
        end
        33962:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        33963:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        33964:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        33965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        33999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34088:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd36;
        end
        34089:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd218;
        end
        34090:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34091:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd146;
        end
        34092:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        34093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34096:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        34097:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34098:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        34099:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        34100:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34101:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        34102:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd18;
        end
        34103:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd195;
        end
        34104:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34105:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd134;
        end
        34106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd21;
        end
        34107:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd123;
        end
        34108:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd0;
        end
        34109:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        34110:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34111:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34112:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34113:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd109;
        end
        34114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34119:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        34120:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34121:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd183;
        end
        34122:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd163;
        end
        34123:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34124:
        begin
            RED=8'd0;
            GRN=8'd122;
            BLU=8'd145;
        end
        34125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34126:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd146;
        end
        34127:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34128:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd193;
        end
        34129:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd105;
        end
        34130:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34131:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd166;
        end
        34132:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd183;
        end
        34133:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34134:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34135:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd147;
        end
        34136:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd5;
        end
        34137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd23;
        end
        34138:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd208;
        end
        34139:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34140:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd112;
        end
        34141:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd186;
        end
        34142:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34143:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd77;
        end
        34144:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        34145:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34146:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        34147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34151:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        34152:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        34153:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34154:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        34155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd35;
        end
        34156:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd227;
        end
        34157:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34158:
        begin
            RED=8'd0;
            GRN=8'd79;
            BLU=8'd88;
        end
        34159:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd195;
        end
        34160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34161:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd156;
        end
        34162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34166:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        34167:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34168:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34169:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34170:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34171:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd227;
        end
        34172:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd49;
        end
        34173:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        34174:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34175:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        34176:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd0;
        end
        34177:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd18;
        end
        34178:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd43;
        end
        34179:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd212;
        end
        34180:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34181:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd212;
        end
        34182:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd28;
        end
        34183:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd207;
        end
        34184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34185:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd151;
        end
        34186:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd180;
        end
        34187:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd86;
        end
        34188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34192:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd91;
        end
        34193:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd198;
        end
        34194:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd95;
        end
        34195:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        34196:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34197:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd41;
        end
        34198:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd91;
        end
        34199:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34200:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd220;
        end
        34201:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd89;
        end
        34202:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd232;
        end
        34203:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34204:
        begin
            RED=8'd0;
            GRN=8'd66;
            BLU=8'd56;
        end
        34205:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd5;
        end
        34206:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd38;
        end
        34207:
        begin
            RED=8'd0;
            GRN=8'd97;
            BLU=8'd170;
        end
        34208:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34210:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd68;
        end
        34211:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        34212:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34213:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        34214:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        34215:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        34216:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34217:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd129;
        end
        34218:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        34219:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34220:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        34221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34344:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd36;
        end
        34345:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd218;
        end
        34346:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34347:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd146;
        end
        34348:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        34349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34352:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        34353:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34354:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        34355:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        34356:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34357:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        34358:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd23;
        end
        34359:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd204;
        end
        34360:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34361:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd134;
        end
        34362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        34363:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd7;
        end
        34364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34365:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        34366:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34367:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34368:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34369:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd150;
        end
        34370:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        34371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34375:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        34376:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34377:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        34378:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd90;
        end
        34379:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34380:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd210;
        end
        34381:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd26;
        end
        34382:
        begin
            RED=8'd0;
            GRN=8'd90;
            BLU=8'd161;
        end
        34383:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34384:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd230;
        end
        34385:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd225;
        end
        34386:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34387:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd174;
        end
        34388:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd152;
        end
        34389:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34390:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34391:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd227;
        end
        34392:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd86;
        end
        34393:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd31;
        end
        34394:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd215;
        end
        34395:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34396:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd225;
        end
        34397:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd229;
        end
        34398:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34399:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd92;
        end
        34400:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        34401:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34402:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        34403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34407:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        34408:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        34409:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34410:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        34411:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd48;
        end
        34412:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        34413:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34414:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd86;
        end
        34415:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd183;
        end
        34416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34417:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd156;
        end
        34418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34422:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        34423:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34424:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34425:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34426:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd220;
        end
        34427:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd113;
        end
        34428:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd3;
        end
        34429:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        34430:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34431:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        34432:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd0;
        end
        34433:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd32;
        end
        34434:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd201;
        end
        34435:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd231;
        end
        34436:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34437:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd212;
        end
        34438:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd28;
        end
        34439:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd179;
        end
        34440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34441:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd200;
        end
        34442:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd218;
        end
        34443:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd49;
        end
        34444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34448:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd128;
        end
        34449:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd171;
        end
        34450:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd65;
        end
        34451:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd229;
        end
        34452:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34453:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd78;
        end
        34454:
        begin
            RED=8'd0;
            GRN=8'd27;
            BLU=8'd77;
        end
        34455:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34456:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd223;
        end
        34457:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd101;
        end
        34458:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd232;
        end
        34459:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd221;
        end
        34460:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd41;
        end
        34461:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd9;
        end
        34462:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd167;
        end
        34463:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd228;
        end
        34464:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34465:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34466:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd68;
        end
        34467:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        34468:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34469:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        34470:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        34471:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        34472:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34473:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd116;
        end
        34474:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        34475:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34476:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        34477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34600:
        begin
            RED=8'd0;
            GRN=8'd10;
            BLU=8'd36;
        end
        34601:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd218;
        end
        34602:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34603:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd146;
        end
        34604:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        34605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34606:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd163;
        end
        34607:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd83;
        end
        34608:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        34609:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34610:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        34611:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        34612:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34613:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        34614:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd23;
        end
        34615:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd205;
        end
        34616:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34617:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd134;
        end
        34618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34621:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        34622:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34623:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34624:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34625:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd180;
        end
        34626:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd6;
        end
        34627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34631:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        34632:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34633:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        34634:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd71;
        end
        34635:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        34636:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd226;
        end
        34637:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd54;
        end
        34638:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd162;
        end
        34639:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34640:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd198;
        end
        34641:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd35;
        end
        34642:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd31;
        end
        34643:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd24;
        end
        34644:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd100;
        end
        34645:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34646:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34647:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34648:
        begin
            RED=8'd0;
            GRN=8'd146;
            BLU=8'd186;
        end
        34649:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd32;
        end
        34650:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd215;
        end
        34651:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34652:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd128;
        end
        34653:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd31;
        end
        34654:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd31;
        end
        34655:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd14;
        end
        34656:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        34657:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34658:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        34659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34663:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        34664:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        34665:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34666:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        34667:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd49;
        end
        34668:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        34669:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34670:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd86;
        end
        34671:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd182;
        end
        34672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34673:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd169;
        end
        34674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34678:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        34679:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34680:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd225;
        end
        34681:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd69;
        end
        34682:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd30;
        end
        34683:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd14;
        end
        34684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34685:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        34686:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34687:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        34688:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd15;
        end
        34689:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd177;
        end
        34690:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd226;
        end
        34691:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd173;
        end
        34692:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34693:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd212;
        end
        34694:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd28;
        end
        34695:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd150;
        end
        34696:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34697:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        34698:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd211;
        end
        34699:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd30;
        end
        34700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34704:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd156;
        end
        34705:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd144;
        end
        34706:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd44;
        end
        34707:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd223;
        end
        34708:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34709:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd106;
        end
        34710:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd34;
        end
        34711:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd217;
        end
        34712:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd228;
        end
        34713:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd169;
        end
        34714:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        34715:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd172;
        end
        34716:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd5;
        end
        34717:
        begin
            RED=8'd0;
            GRN=8'd64;
            BLU=8'd138;
        end
        34718:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd224;
        end
        34719:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd170;
        end
        34720:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34721:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34722:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd68;
        end
        34723:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        34724:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34725:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        34726:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        34727:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        34728:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34729:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd116;
        end
        34730:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        34731:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34732:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        34733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34856:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd19;
        end
        34857:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd209;
        end
        34858:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34859:
        begin
            RED=8'd0;
            GRN=8'd134;
            BLU=8'd162;
        end
        34860:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd2;
        end
        34861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34862:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd178;
        end
        34863:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd119;
        end
        34864:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        34865:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34866:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        34867:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        34868:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34869:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        34870:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd23;
        end
        34871:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd205;
        end
        34872:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34873:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd134;
        end
        34874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34875:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd124;
        end
        34876:
        begin
            RED=8'd0;
            GRN=8'd35;
            BLU=8'd42;
        end
        34877:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        34878:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34879:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34880:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34881:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd213;
        end
        34882:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd12;
        end
        34883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34887:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        34888:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34889:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        34890:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd69;
        end
        34891:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        34892:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        34893:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd65;
        end
        34894:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd162;
        end
        34895:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34896:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd193;
        end
        34897:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd4;
        end
        34898:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd39;
        end
        34899:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd8;
        end
        34900:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd29;
        end
        34901:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd195;
        end
        34902:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34903:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34904:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd221;
        end
        34905:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd76;
        end
        34906:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd215;
        end
        34907:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34908:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd112;
        end
        34909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        34910:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd44;
        end
        34911:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd2;
        end
        34912:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        34913:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34914:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        34915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34919:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        34920:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        34921:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34922:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        34923:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd49;
        end
        34924:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd228;
        end
        34925:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34926:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd86;
        end
        34927:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd182;
        end
        34928:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34929:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd159;
        end
        34930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34934:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        34935:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34936:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        34937:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        34938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34941:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        34942:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34943:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        34944:
        begin
            RED=8'd0;
            GRN=8'd34;
            BLU=8'd54;
        end
        34945:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd225;
        end
        34946:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd216;
        end
        34947:
        begin
            RED=8'd0;
            GRN=8'd81;
            BLU=8'd129;
        end
        34948:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34949:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd212;
        end
        34950:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd28;
        end
        34951:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd108;
        end
        34952:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34953:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34954:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd197;
        end
        34955:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd14;
        end
        34956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34960:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd172;
        end
        34961:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd212;
        end
        34962:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd191;
        end
        34963:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd230;
        end
        34964:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34965:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd121;
        end
        34966:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd6;
        end
        34967:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd149;
        end
        34968:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd231;
        end
        34969:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd220;
        end
        34970:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd221;
        end
        34971:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd65;
        end
        34972:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd14;
        end
        34973:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd206;
        end
        34974:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34975:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd112;
        end
        34976:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34977:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34978:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd68;
        end
        34979:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        34980:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34981:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        34982:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        34983:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        34984:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34985:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd116;
        end
        34986:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        34987:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        34988:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        34989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        34999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        35113:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd202;
        end
        35114:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35115:
        begin
            RED=8'd0;
            GRN=8'd142;
            BLU=8'd176;
        end
        35116:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd3;
        end
        35117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35118:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd186;
        end
        35119:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd125;
        end
        35120:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        35121:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35122:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        35123:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        35124:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35125:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        35126:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd23;
        end
        35127:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd205;
        end
        35128:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35129:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd134;
        end
        35130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35131:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd168;
        end
        35132:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd95;
        end
        35133:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        35134:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35135:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35136:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35137:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd229;
        end
        35138:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd31;
        end
        35139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35143:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        35144:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35145:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        35146:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd69;
        end
        35147:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd232;
        end
        35148:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35149:
        begin
            RED=8'd0;
            GRN=8'd82;
            BLU=8'd82;
        end
        35150:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd162;
        end
        35151:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35152:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd193;
        end
        35153:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd4;
        end
        35154:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd103;
        end
        35155:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd126;
        end
        35156:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd52;
        end
        35157:
        begin
            RED=8'd0;
            GRN=8'd82;
            BLU=8'd125;
        end
        35158:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd221;
        end
        35159:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35160:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        35161:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd104;
        end
        35162:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd215;
        end
        35163:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35164:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd112;
        end
        35165:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd10;
        end
        35166:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd156;
        end
        35167:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd66;
        end
        35168:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        35169:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35170:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        35171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35175:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        35176:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        35177:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35178:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        35179:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd39;
        end
        35180:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd227;
        end
        35181:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35182:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd87;
        end
        35183:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd191;
        end
        35184:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35185:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd156;
        end
        35186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35190:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        35191:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35192:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        35193:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        35194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35197:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        35198:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35199:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        35200:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd98;
        end
        35201:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        35202:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd209;
        end
        35203:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd108;
        end
        35204:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35205:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd212;
        end
        35206:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd28;
        end
        35207:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd76;
        end
        35208:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35209:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35210:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd166;
        end
        35211:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd3;
        end
        35212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd8;
        end
        35216:
        begin
            RED=8'd0;
            GRN=8'd116;
            BLU=8'd191;
        end
        35217:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35218:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35219:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35220:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35221:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd148;
        end
        35222:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd6;
        end
        35223:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd160;
        end
        35224:
        begin
            RED=8'd0;
            GRN=8'd140;
            BLU=8'd180;
        end
        35225:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd81;
        end
        35226:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd65;
        end
        35227:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd11;
        end
        35228:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd45;
        end
        35229:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd224;
        end
        35230:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35231:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd84;
        end
        35232:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35233:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35234:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd68;
        end
        35235:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        35236:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35237:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        35238:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        35239:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        35240:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35241:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd116;
        end
        35242:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        35243:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35244:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        35245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35369:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd174;
        end
        35370:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35371:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd189;
        end
        35372:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd5;
        end
        35373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35374:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd198;
        end
        35375:
        begin
            RED=8'd0;
            GRN=8'd95;
            BLU=8'd101;
        end
        35376:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        35377:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35378:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        35379:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        35380:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35381:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        35382:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd16;
        end
        35383:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd192;
        end
        35384:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35385:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd143;
        end
        35386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35387:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd182;
        end
        35388:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd103;
        end
        35389:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        35390:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35391:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd224;
        end
        35392:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35393:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35394:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd67;
        end
        35395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35399:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        35400:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35401:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        35402:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd55;
        end
        35403:
        begin
            RED=8'd0;
            GRN=8'd154;
            BLU=8'd232;
        end
        35404:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35405:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd89;
        end
        35406:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd141;
        end
        35407:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35408:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd201;
        end
        35409:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd5;
        end
        35410:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd126;
        end
        35411:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd161;
        end
        35412:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd156;
        end
        35413:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd107;
        end
        35414:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd128;
        end
        35415:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd232;
        end
        35416:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35417:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd99;
        end
        35418:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd206;
        end
        35419:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35420:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd121;
        end
        35421:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd12;
        end
        35422:
        begin
            RED=8'd0;
            GRN=8'd121;
            BLU=8'd199;
        end
        35423:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd72;
        end
        35424:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        35425:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35426:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        35427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35431:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd23;
        end
        35432:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd222;
        end
        35433:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35434:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        35435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd25;
        end
        35436:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd226;
        end
        35437:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35438:
        begin
            RED=8'd0;
            GRN=8'd84;
            BLU=8'd97;
        end
        35439:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd195;
        end
        35440:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35441:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd136;
        end
        35442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35446:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        35447:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35448:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        35449:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        35450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35453:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        35454:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35455:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        35456:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd121;
        end
        35457:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35458:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd211;
        end
        35459:
        begin
            RED=8'd0;
            GRN=8'd79;
            BLU=8'd122;
        end
        35460:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35461:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd212;
        end
        35462:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd28;
        end
        35463:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd43;
        end
        35464:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd232;
        end
        35465:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35466:
        begin
            RED=8'd0;
            GRN=8'd116;
            BLU=8'd136;
        end
        35467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35471:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd23;
        end
        35472:
        begin
            RED=8'd0;
            GRN=8'd132;
            BLU=8'd207;
        end
        35473:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd124;
        end
        35474:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd88;
        end
        35475:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd210;
        end
        35476:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35477:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd178;
        end
        35478:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd41;
        end
        35479:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd209;
        end
        35480:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd124;
        end
        35481:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd6;
        end
        35482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35484:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd64;
        end
        35485:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd229;
        end
        35486:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35487:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd101;
        end
        35488:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35489:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35490:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd68;
        end
        35491:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        35492:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35493:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        35494:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        35495:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        35496:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35497:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd116;
        end
        35498:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        35499:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35500:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        35501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35625:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd121;
        end
        35626:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35627:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd214;
        end
        35628:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd9;
        end
        35629:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd21;
        end
        35630:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd209;
        end
        35631:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd65;
        end
        35632:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        35633:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35634:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        35635:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        35636:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35637:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        35638:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd8;
        end
        35639:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd162;
        end
        35640:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35641:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd156;
        end
        35642:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        35643:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd196;
        end
        35644:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd76;
        end
        35645:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        35646:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35647:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd166;
        end
        35648:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd232;
        end
        35649:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35650:
        begin
            RED=8'd0;
            GRN=8'd94;
            BLU=8'd100;
        end
        35651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35655:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        35656:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35657:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        35658:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd47;
        end
        35659:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd232;
        end
        35660:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35661:
        begin
            RED=8'd0;
            GRN=8'd90;
            BLU=8'd98;
        end
        35662:
        begin
            RED=8'd0;
            GRN=8'd49;
            BLU=8'd102;
        end
        35663:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35664:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd220;
        end
        35665:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd6;
        end
        35666:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd134;
        end
        35667:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd133;
        end
        35668:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd202;
        end
        35669:
        begin
            RED=8'd0;
            GRN=8'd111;
            BLU=8'd126;
        end
        35670:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd42;
        end
        35671:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd212;
        end
        35672:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd229;
        end
        35673:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd73;
        end
        35674:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd181;
        end
        35675:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35676:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd141;
        end
        35677:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd14;
        end
        35678:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd200;
        end
        35679:
        begin
            RED=8'd0;
            GRN=8'd52;
            BLU=8'd45;
        end
        35680:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd211;
        end
        35681:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35682:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd112;
        end
        35683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35687:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd21;
        end
        35688:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd217;
        end
        35689:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35690:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd87;
        end
        35691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd9;
        end
        35692:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd209;
        end
        35693:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35694:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd113;
        end
        35695:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd208;
        end
        35696:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35697:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd97;
        end
        35698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35702:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        35703:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35704:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        35705:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        35706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35709:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        35710:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35711:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        35712:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd118;
        end
        35713:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35714:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd217;
        end
        35715:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd163;
        end
        35716:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35717:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd212;
        end
        35718:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd28;
        end
        35719:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd21;
        end
        35720:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd216;
        end
        35721:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        35722:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd98;
        end
        35723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35727:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd38;
        end
        35728:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd220;
        end
        35729:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd42;
        end
        35730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35731:
        begin
            RED=8'd0;
            GRN=8'd104;
            BLU=8'd180;
        end
        35732:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35733:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd198;
        end
        35734:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd86;
        end
        35735:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd232;
        end
        35736:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd173;
        end
        35737:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd125;
        end
        35738:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd125;
        end
        35739:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd105;
        end
        35740:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd74;
        end
        35741:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd228;
        end
        35742:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35743:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd148;
        end
        35744:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35745:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35746:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd68;
        end
        35747:
        begin
            RED=8'd0;
            GRN=8'd93;
            BLU=8'd161;
        end
        35748:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35749:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        35750:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        35751:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        35752:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35753:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd116;
        end
        35754:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        35755:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35756:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        35757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35881:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd51;
        end
        35882:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd220;
        end
        35883:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35884:
        begin
            RED=8'd0;
            GRN=8'd67;
            BLU=8'd62;
        end
        35885:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd90;
        end
        35886:
        begin
            RED=8'd0;
            GRN=8'd145;
            BLU=8'd198;
        end
        35887:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd26;
        end
        35888:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        35889:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35890:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        35891:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        35892:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35893:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        35894:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd4;
        end
        35895:
        begin
            RED=8'd0;
            GRN=8'd56;
            BLU=8'd107;
        end
        35896:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd230;
        end
        35897:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd183;
        end
        35898:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd28;
        end
        35899:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd208;
        end
        35900:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd47;
        end
        35901:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        35902:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35903:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd122;
        end
        35904:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd219;
        end
        35905:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35906:
        begin
            RED=8'd0;
            GRN=8'd120;
            BLU=8'd138;
        end
        35907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35911:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        35912:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35913:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        35914:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd47;
        end
        35915:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd232;
        end
        35916:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35917:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd113;
        end
        35918:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd48;
        end
        35919:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd226;
        end
        35920:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35921:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd51;
        end
        35922:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd165;
        end
        35923:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd84;
        end
        35924:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd169;
        end
        35925:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd176;
        end
        35926:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd38;
        end
        35927:
        begin
            RED=8'd0;
            GRN=8'd128;
            BLU=8'd205;
        end
        35928:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd221;
        end
        35929:
        begin
            RED=8'd0;
            GRN=8'd40;
            BLU=8'd30;
        end
        35930:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd127;
        end
        35931:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35932:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd185;
        end
        35933:
        begin
            RED=8'd0;
            GRN=8'd32;
            BLU=8'd42;
        end
        35934:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd194;
        end
        35935:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd22;
        end
        35936:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd199;
        end
        35937:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35938:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd167;
        end
        35939:
        begin
            RED=8'd0;
            GRN=8'd45;
            BLU=8'd51;
        end
        35940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35943:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd17;
        end
        35944:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd207;
        end
        35945:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35946:
        begin
            RED=8'd0;
            GRN=8'd122;
            BLU=8'd154;
        end
        35947:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd40;
        end
        35948:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd158;
        end
        35949:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35950:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd145;
        end
        35951:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd225;
        end
        35952:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd226;
        end
        35953:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd43;
        end
        35954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35958:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        35959:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35960:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        35961:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        35962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35965:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        35966:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35967:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        35968:
        begin
            RED=8'd0;
            GRN=8'd57;
            BLU=8'd90;
        end
        35969:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        35970:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd226;
        end
        35971:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd208;
        end
        35972:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35973:
        begin
            RED=8'd0;
            GRN=8'd159;
            BLU=8'd221;
        end
        35974:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd77;
        end
        35975:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd11;
        end
        35976:
        begin
            RED=8'd0;
            GRN=8'd116;
            BLU=8'd191;
        end
        35977:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd230;
        end
        35978:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd63;
        end
        35979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35983:
        begin
            RED=8'd0;
            GRN=8'd23;
            BLU=8'd48;
        end
        35984:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd229;
        end
        35985:
        begin
            RED=8'd0;
            GRN=8'd36;
            BLU=8'd17;
        end
        35986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        35987:
        begin
            RED=8'd0;
            GRN=8'd82;
            BLU=8'd152;
        end
        35988:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35989:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd217;
        end
        35990:
        begin
            RED=8'd0;
            GRN=8'd71;
            BLU=8'd114;
        end
        35991:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35992:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35993:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35994:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35995:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd211;
        end
        35996:
        begin
            RED=8'd0;
            GRN=8'd76;
            BLU=8'd108;
        end
        35997:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd223;
        end
        35998:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        35999:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd202;
        end
        36000:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36001:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36002:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd125;
        end
        36003:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd161;
        end
        36004:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36005:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        36006:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        36007:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        36008:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36009:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd116;
        end
        36010:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        36011:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36012:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        36013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36137:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        36138:
        begin
            RED=8'd0;
            GRN=8'd97;
            BLU=8'd149;
        end
        36139:
        begin
            RED=8'd0;
            GRN=8'd152;
            BLU=8'd221;
        end
        36140:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd164;
        end
        36141:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd166;
        end
        36142:
        begin
            RED=8'd0;
            GRN=8'd101;
            BLU=8'd126;
        end
        36143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36144:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd185;
        end
        36145:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36146:
        begin
            RED=8'd0;
            GRN=8'd124;
            BLU=8'd148;
        end
        36147:
        begin
            RED=8'd0;
            GRN=8'd62;
            BLU=8'd110;
        end
        36148:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36149:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd219;
        end
        36150:
        begin
            RED=8'd0;
            GRN=8'd19;
            BLU=8'd4;
        end
        36151:
        begin
            RED=8'd0;
            GRN=8'd18;
            BLU=8'd40;
        end
        36152:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd194;
        end
        36153:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd216;
        end
        36154:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd126;
        end
        36155:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd168;
        end
        36156:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd21;
        end
        36157:
        begin
            RED=8'd0;
            GRN=8'd129;
            BLU=8'd213;
        end
        36158:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36159:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd122;
        end
        36160:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd187;
        end
        36161:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36162:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd178;
        end
        36163:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd0;
        end
        36164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36167:
        begin
            RED=8'd0;
            GRN=8'd123;
            BLU=8'd206;
        end
        36168:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36169:
        begin
            RED=8'd0;
            GRN=8'd147;
            BLU=8'd182;
        end
        36170:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd42;
        end
        36171:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd226;
        end
        36172:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36173:
        begin
            RED=8'd0;
            GRN=8'd113;
            BLU=8'd132;
        end
        36174:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd6;
        end
        36175:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd168;
        end
        36176:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd230;
        end
        36177:
        begin
            RED=8'd0;
            GRN=8'd119;
            BLU=8'd152;
        end
        36178:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd177;
        end
        36179:
        begin
            RED=8'd0;
            GRN=8'd37;
            BLU=8'd31;
        end
        36180:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd93;
        end
        36181:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd209;
        end
        36182:
        begin
            RED=8'd0;
            GRN=8'd92;
            BLU=8'd129;
        end
        36183:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd218;
        end
        36184:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd161;
        end
        36185:
        begin
            RED=8'd0;
            GRN=8'd14;
            BLU=8'd0;
        end
        36186:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd52;
        end
        36187:
        begin
            RED=8'd0;
            GRN=8'd133;
            BLU=8'd205;
        end
        36188:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd225;
        end
        36189:
        begin
            RED=8'd0;
            GRN=8'd97;
            BLU=8'd132;
        end
        36190:
        begin
            RED=8'd0;
            GRN=8'd117;
            BLU=8'd144;
        end
        36191:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd6;
        end
        36192:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd155;
        end
        36193:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd232;
        end
        36194:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd221;
        end
        36195:
        begin
            RED=8'd0;
            GRN=8'd75;
            BLU=8'd80;
        end
        36196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36199:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd9;
        end
        36200:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd170;
        end
        36201:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        36202:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd216;
        end
        36203:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd61;
        end
        36204:
        begin
            RED=8'd0;
            GRN=8'd38;
            BLU=8'd75;
        end
        36205:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd212;
        end
        36206:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd196;
        end
        36207:
        begin
            RED=8'd0;
            GRN=8'd155;
            BLU=8'd229;
        end
        36208:
        begin
            RED=8'd0;
            GRN=8'd125;
            BLU=8'd166;
        end
        36209:
        begin
            RED=8'd0;
            GRN=8'd12;
            BLU=8'd3;
        end
        36210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36214:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd120;
        end
        36215:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36216:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd224;
        end
        36217:
        begin
            RED=8'd0;
            GRN=8'd47;
            BLU=8'd44;
        end
        36218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36221:
        begin
            RED=8'd0;
            GRN=8'd63;
            BLU=8'd118;
        end
        36222:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36223:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd215;
        end
        36224:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd44;
        end
        36225:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd211;
        end
        36226:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36227:
        begin
            RED=8'd0;
            GRN=8'd148;
            BLU=8'd211;
        end
        36228:
        begin
            RED=8'd0;
            GRN=8'd153;
            BLU=8'd226;
        end
        36229:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36230:
        begin
            RED=8'd0;
            GRN=8'd126;
            BLU=8'd141;
        end
        36231:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd5;
        end
        36232:
        begin
            RED=8'd0;
            GRN=8'd97;
            BLU=8'd168;
        end
        36233:
        begin
            RED=8'd0;
            GRN=8'd160;
            BLU=8'd226;
        end
        36234:
        begin
            RED=8'd0;
            GRN=8'd41;
            BLU=8'd30;
        end
        36235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36239:
        begin
            RED=8'd0;
            GRN=8'd30;
            BLU=8'd67;
        end
        36240:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd222;
        end
        36241:
        begin
            RED=8'd0;
            GRN=8'd20;
            BLU=8'd5;
        end
        36242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36243:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd126;
        end
        36244:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36245:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36246:
        begin
            RED=8'd0;
            GRN=8'd83;
            BLU=8'd111;
        end
        36247:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd229;
        end
        36248:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36249:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36250:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36251:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36252:
        begin
            RED=8'd0;
            GRN=8'd118;
            BLU=8'd153;
        end
        36253:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd186;
        end
        36254:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36255:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd221;
        end
        36256:
        begin
            RED=8'd0;
            GRN=8'd144;
            BLU=8'd217;
        end
        36257:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36258:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd195;
        end
        36259:
        begin
            RED=8'd0;
            GRN=8'd116;
            BLU=8'd167;
        end
        36260:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36261:
        begin
            RED=8'd0;
            GRN=8'd137;
            BLU=8'd172;
        end
        36262:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        36263:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd222;
        end
        36264:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36265:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd116;
        end
        36266:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd181;
        end
        36267:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36268:
        begin
            RED=8'd0;
            GRN=8'd130;
            BLU=8'd158;
        end
        36269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36394:
        begin
            RED=8'd0;
            GRN=8'd24;
            BLU=8'd39;
        end
        36395:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd143;
        end
        36396:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36397:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd133;
        end
        36398:
        begin
            RED=8'd0;
            GRN=8'd21;
            BLU=8'd27;
        end
        36399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36400:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd130;
        end
        36401:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36402:
        begin
            RED=8'd0;
            GRN=8'd87;
            BLU=8'd104;
        end
        36403:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd77;
        end
        36404:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36405:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd154;
        end
        36406:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd3;
        end
        36407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36408:
        begin
            RED=8'd0;
            GRN=8'd53;
            BLU=8'd97;
        end
        36409:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36410:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36411:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd65;
        end
        36412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36413:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd150;
        end
        36414:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36415:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd85;
        end
        36416:
        begin
            RED=8'd0;
            GRN=8'd60;
            BLU=8'd112;
        end
        36417:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36418:
        begin
            RED=8'd0;
            GRN=8'd105;
            BLU=8'd138;
        end
        36419:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd0;
        end
        36420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36423:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd145;
        end
        36424:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36425:
        begin
            RED=8'd0;
            GRN=8'd103;
            BLU=8'd128;
        end
        36426:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd24;
        end
        36427:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd153;
        end
        36428:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36429:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd105;
        end
        36430:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        36431:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd58;
        end
        36432:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd159;
        end
        36433:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36434:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd105;
        end
        36435:
        begin
            RED=8'd0;
            GRN=8'd5;
            BLU=8'd4;
        end
        36436:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd15;
        end
        36437:
        begin
            RED=8'd0;
            GRN=8'd78;
            BLU=8'd136;
        end
        36438:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36439:
        begin
            RED=8'd0;
            GRN=8'd109;
            BLU=8'd156;
        end
        36440:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd51;
        end
        36441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36443:
        begin
            RED=8'd0;
            GRN=8'd61;
            BLU=8'd112;
        end
        36444:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd163;
        end
        36445:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd159;
        end
        36446:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd53;
        end
        36447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36448:
        begin
            RED=8'd0;
            GRN=8'd28;
            BLU=8'd67;
        end
        36449:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd163;
        end
        36450:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd143;
        end
        36451:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd20;
        end
        36452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36456:
        begin
            RED=8'd0;
            GRN=8'd39;
            BLU=8'd84;
        end
        36457:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd163;
        end
        36458:
        begin
            RED=8'd0;
            GRN=8'd107;
            BLU=8'd134;
        end
        36459:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd13;
        end
        36460:
        begin
            RED=8'd0;
            GRN=8'd4;
            BLU=8'd8;
        end
        36461:
        begin
            RED=8'd0;
            GRN=8'd70;
            BLU=8'd126;
        end
        36462:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd163;
        end
        36463:
        begin
            RED=8'd0;
            GRN=8'd110;
            BLU=8'd158;
        end
        36464:
        begin
            RED=8'd0;
            GRN=8'd46;
            BLU=8'd54;
        end
        36465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36470:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd84;
        end
        36471:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36472:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd157;
        end
        36473:
        begin
            RED=8'd0;
            GRN=8'd33;
            BLU=8'd31;
        end
        36474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36477:
        begin
            RED=8'd0;
            GRN=8'd44;
            BLU=8'd83;
        end
        36478:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36479:
        begin
            RED=8'd0;
            GRN=8'd112;
            BLU=8'd151;
        end
        36480:
        begin
            RED=8'd0;
            GRN=8'd11;
            BLU=8'd7;
        end
        36481:
        begin
            RED=8'd0;
            GRN=8'd74;
            BLU=8'd124;
        end
        36482:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36483:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd124;
        end
        36484:
        begin
            RED=8'd0;
            GRN=8'd98;
            BLU=8'd153;
        end
        36485:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36486:
        begin
            RED=8'd0;
            GRN=8'd89;
            BLU=8'd108;
        end
        36487:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd2;
        end
        36488:
        begin
            RED=8'd0;
            GRN=8'd73;
            BLU=8'd137;
        end
        36489:
        begin
            RED=8'd0;
            GRN=8'd157;
            BLU=8'd214;
        end
        36490:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd0;
        end
        36491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36495:
        begin
            RED=8'd0;
            GRN=8'd25;
            BLU=8'd64;
        end
        36496:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd145;
        end
        36497:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd3;
        end
        36498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36499:
        begin
            RED=8'd0;
            GRN=8'd42;
            BLU=8'd79;
        end
        36500:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36501:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36502:
        begin
            RED=8'd0;
            GRN=8'd48;
            BLU=8'd68;
        end
        36503:
        begin
            RED=8'd0;
            GRN=8'd136;
            BLU=8'd209;
        end
        36504:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36505:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36506:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36507:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36508:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd170;
        end
        36509:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd93;
        end
        36510:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36511:
        begin
            RED=8'd0;
            GRN=8'd106;
            BLU=8'd143;
        end
        36512:
        begin
            RED=8'd0;
            GRN=8'd80;
            BLU=8'd135;
        end
        36513:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36514:
        begin
            RED=8'd0;
            GRN=8'd102;
            BLU=8'd140;
        end
        36515:
        begin
            RED=8'd0;
            GRN=8'd85;
            BLU=8'd124;
        end
        36516:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36517:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd121;
        end
        36518:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd0;
        end
        36519:
        begin
            RED=8'd0;
            GRN=8'd96;
            BLU=8'd156;
        end
        36520:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36521:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd82;
        end
        36522:
        begin
            RED=8'd0;
            GRN=8'd72;
            BLU=8'd127;
        end
        36523:
        begin
            RED=8'd0;
            GRN=8'd114;
            BLU=8'd163;
        end
        36524:
        begin
            RED=8'd0;
            GRN=8'd91;
            BLU=8'd111;
        end
        36525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36744:
        begin
            RED=8'd0;
            GRN=8'd50;
            BLU=8'd109;
        end
        36745:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd188;
        end
        36746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36758:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd23;
        end
        36759:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd186;
        end
        36760:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd209;
        end
        36761:
        begin
            RED=8'd0;
            GRN=8'd127;
            BLU=8'd182;
        end
        36762:
        begin
            RED=8'd0;
            GRN=8'd143;
            BLU=8'd211;
        end
        36763:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        36764:
        begin
            RED=8'd0;
            GRN=8'd138;
            BLU=8'd170;
        end
        36765:
        begin
            RED=8'd0;
            GRN=8'd7;
            BLU=8'd4;
        end
        36766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        36998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd3;
        end
        36999:
        begin
            RED=8'd0;
            GRN=8'd13;
            BLU=8'd17;
        end
        37000:
        begin
            RED=8'd0;
            GRN=8'd65;
            BLU=8'd125;
        end
        37001:
        begin
            RED=8'd0;
            GRN=8'd131;
            BLU=8'd157;
        end
        37002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37014:
        begin
            RED=8'd0;
            GRN=8'd29;
            BLU=8'd80;
        end
        37015:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        37016:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd114;
        end
        37017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37018:
        begin
            RED=8'd0;
            GRN=8'd68;
            BLU=8'd127;
        end
        37019:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd232;
        end
        37020:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd166;
        end
        37021:
        begin
            RED=8'd0;
            GRN=8'd6;
            BLU=8'd3;
        end
        37022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37254:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd22;
        end
        37255:
        begin
            RED=8'd0;
            GRN=8'd99;
            BLU=8'd131;
        end
        37256:
        begin
            RED=8'd0;
            GRN=8'd88;
            BLU=8'd153;
        end
        37257:
        begin
            RED=8'd0;
            GRN=8'd100;
            BLU=8'd109;
        end
        37258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37270:
        begin
            RED=8'd0;
            GRN=8'd51;
            BLU=8'd104;
        end
        37271:
        begin
            RED=8'd0;
            GRN=8'd161;
            BLU=8'd232;
        end
        37272:
        begin
            RED=8'd0;
            GRN=8'd55;
            BLU=8'd46;
        end
        37273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        37274:
        begin
            RED=8'd0;
            GRN=8'd31;
            BLU=8'd75;
        end
        37275:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd231;
        end
        37276:
        begin
            RED=8'd0;
            GRN=8'd115;
            BLU=8'd134;
        end
        37277:
        begin
            RED=8'd0;
            GRN=8'd3;
            BLU=8'd0;
        end
        37278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37510:
        begin
            RED=8'd0;
            GRN=8'd43;
            BLU=8'd85;
        end
        37511:
        begin
            RED=8'd0;
            GRN=8'd151;
            BLU=8'd220;
        end
        37512:
        begin
            RED=8'd0;
            GRN=8'd141;
            BLU=8'd202;
        end
        37513:
        begin
            RED=8'd0;
            GRN=8'd58;
            BLU=8'd51;
        end
        37514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37526:
        begin
            RED=8'd0;
            GRN=8'd22;
            BLU=8'd76;
        end
        37527:
        begin
            RED=8'd0;
            GRN=8'd156;
            BLU=8'd232;
        end
        37528:
        begin
            RED=8'd0;
            GRN=8'd108;
            BLU=8'd125;
        end
        37529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd13;
        end
        37530:
        begin
            RED=8'd0;
            GRN=8'd95;
            BLU=8'd160;
        end
        37531:
        begin
            RED=8'd0;
            GRN=8'd162;
            BLU=8'd226;
        end
        37532:
        begin
            RED=8'd0;
            GRN=8'd54;
            BLU=8'd48;
        end
        37533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37766:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd21;
        end
        37767:
        begin
            RED=8'd0;
            GRN=8'd135;
            BLU=8'd210;
        end
        37768:
        begin
            RED=8'd0;
            GRN=8'd149;
            BLU=8'd192;
        end
        37769:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd13;
        end
        37770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37782:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd10;
        end
        37783:
        begin
            RED=8'd0;
            GRN=8'd86;
            BLU=8'd150;
        end
        37784:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd226;
        end
        37785:
        begin
            RED=8'd0;
            GRN=8'd158;
            BLU=8'd226;
        end
        37786:
        begin
            RED=8'd0;
            GRN=8'd150;
            BLU=8'd216;
        end
        37787:
        begin
            RED=8'd0;
            GRN=8'd77;
            BLU=8'd79;
        end
        37788:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        37789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        37999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        38023:
        begin
            RED=8'd0;
            GRN=8'd15;
            BLU=8'd23;
        end
        38024:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd21;
        end
        38025:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd1;
        end
        38026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        38039:
        begin
            RED=8'd0;
            GRN=8'd9;
            BLU=8'd16;
        end
        38040:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd25;
        end
        38041:
        begin
            RED=8'd0;
            GRN=8'd17;
            BLU=8'd25;
        end
        38042:
        begin
            RED=8'd0;
            GRN=8'd16;
            BLU=8'd24;
        end
        38043:
        begin
            RED=8'd0;
            GRN=8'd8;
            BLU=8'd8;
        end
        38044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38150:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38151:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38156:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38157:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38158:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38159:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38160:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38161:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38162:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38163:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38164:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38165:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38166:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38167:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38406:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38407:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38408:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38409:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38410:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38411:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38412:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38413:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38414:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38415:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38416:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38417:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38418:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38419:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38420:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38421:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38422:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38423:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38662:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38663:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38664:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38665:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38666:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38667:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38668:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38669:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38670:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38671:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38672:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38673:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38674:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38675:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38676:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38677:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38678:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38679:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        38999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39169:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39172:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39173:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39174:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39175:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39176:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39177:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39178:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39179:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39180:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39181:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39182:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39183:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39184:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39185:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39186:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39187:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39188:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39189:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39190:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39191:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39424:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39425:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39426:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39427:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39428:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39429:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39430:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39431:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39432:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39433:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39434:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39435:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39436:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39437:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39438:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39439:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39440:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39441:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39442:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39443:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39444:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39445:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39446:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39447:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39680:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39681:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39682:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39683:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39684:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39685:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39686:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39687:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39688:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39689:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39690:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39691:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39692:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39693:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39694:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39695:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39696:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39697:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39698:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39699:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39700:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39701:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39702:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39703:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39984:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39985:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39986:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39987:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39988:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39989:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39990:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39991:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        39999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40120:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40121:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40122:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40123:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40124:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40125:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40126:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40127:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40134:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40135:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40136:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40137:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40138:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40139:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40140:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40141:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40142:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40143:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40144:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40146:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40148:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40149:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40192:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40193:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40194:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40195:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40196:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40197:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40198:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40199:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40200:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40201:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40202:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40203:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40204:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40205:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40206:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40207:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40208:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40209:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40210:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40212:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40213:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40214:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40215:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40221:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40222:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40223:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40225:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40226:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40227:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40228:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40229:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40230:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40231:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40236:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40237:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40238:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40239:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40240:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40241:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40248:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40249:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40250:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40251:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40252:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40253:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40254:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40255:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40260:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40261:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40262:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40263:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40264:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40265:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40266:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40267:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40268:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40269:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40270:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40271:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40272:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40273:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40274:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40275:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40276:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40277:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40278:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40279:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40280:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40281:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40282:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40283:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40284:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40285:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40286:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40287:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40288:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40289:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40290:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40291:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40292:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40293:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40294:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40295:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40296:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40297:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40298:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40299:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40300:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40301:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40302:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40303:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40304:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40305:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40306:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40307:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40308:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40309:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40310:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40311:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40312:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40313:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40314:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40315:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40316:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40317:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40318:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40319:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40320:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40321:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40322:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40323:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40324:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40325:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40326:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40327:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40328:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40329:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40330:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40331:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40332:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40333:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40334:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40335:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40336:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40337:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40338:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40339:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40340:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40341:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40342:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40344:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40345:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40346:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40347:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40348:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40349:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40350:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40351:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40354:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40355:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40356:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40357:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40358:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40359:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40360:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40361:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40362:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40363:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40364:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40365:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40366:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40367:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40368:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40369:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40370:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40371:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40376:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40377:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40378:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40379:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40380:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40381:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40382:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40383:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40386:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40387:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40388:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40389:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40390:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40391:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40392:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40393:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40394:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40395:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40396:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40397:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40398:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40399:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40400:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40401:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40402:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40403:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40404:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40405:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40448:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40449:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40450:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40451:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40452:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40453:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40454:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40455:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40456:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40457:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40458:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40459:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40460:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40461:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40462:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40463:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40464:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40465:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40466:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40467:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40468:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40469:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40472:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40473:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40474:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40475:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40476:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40477:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40478:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40479:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40483:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40484:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40485:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40486:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40487:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40488:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40489:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40490:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40491:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40492:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40493:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40494:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40495:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40496:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40497:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40498:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40499:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40500:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40501:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40504:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40505:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40506:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40507:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40508:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40509:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40510:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40511:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40513:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40514:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40515:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40516:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40517:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40518:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40519:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40520:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40521:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40522:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40523:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40524:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40525:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40526:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40527:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40528:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40529:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40530:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40531:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40532:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40533:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40534:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40535:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40536:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40537:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40538:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40539:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40540:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40541:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40542:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40543:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40544:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40545:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40546:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40547:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40548:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40549:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40550:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40551:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40552:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40553:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40554:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40555:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40556:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40557:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40558:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40559:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40560:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40561:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40562:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40563:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40564:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40565:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40566:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40567:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40568:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40569:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40570:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40571:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40572:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40573:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40574:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40575:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40576:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40577:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40578:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40579:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40580:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40581:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40582:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40583:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40584:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40585:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40586:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40587:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40588:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40589:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40590:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40591:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40592:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40593:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40594:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40595:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40596:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40600:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40601:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40602:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40603:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40604:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40605:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40606:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40607:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40614:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40615:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40616:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40617:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40618:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40619:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40620:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40621:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40622:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40623:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40624:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40625:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40626:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40627:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40628:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40629:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40630:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40632:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40633:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40634:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40635:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40636:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40637:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40638:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40639:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40641:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40642:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40643:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40644:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40645:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40646:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40647:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40648:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40649:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40650:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40651:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40652:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40653:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40654:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40655:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40656:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40657:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40658:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40659:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40660:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40661:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40704:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40705:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40706:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40707:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40708:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40709:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40710:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40711:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40712:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40713:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40714:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40715:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40716:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40717:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40718:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40719:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40720:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40721:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40722:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40728:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40729:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40730:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40731:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40732:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40733:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40734:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40735:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40746:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40747:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40748:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40749:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40750:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40751:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40752:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40753:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40754:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40755:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40756:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40757:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40758:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40759:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40760:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40761:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40762:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40763:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40764:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40765:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40766:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40767:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40768:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40769:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40770:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40771:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40772:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40773:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40774:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40775:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40776:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40777:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40778:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40779:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40780:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40781:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40782:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40783:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40784:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40785:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40786:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40787:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40788:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40789:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40790:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40791:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40792:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40793:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40794:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40795:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40796:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40797:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40798:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40799:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40800:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40801:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40802:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40803:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40804:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40805:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40806:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40807:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40808:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40809:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40810:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40811:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40812:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40813:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40814:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40815:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40816:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40817:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40818:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40819:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40820:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40821:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40822:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40823:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40824:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40825:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40826:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40827:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40828:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40829:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40830:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40831:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40832:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40833:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40834:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40835:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40836:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40837:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40838:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40839:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40840:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40841:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40842:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40843:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40844:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40845:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40856:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40857:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40858:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40859:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40860:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40861:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40862:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40863:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40874:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40875:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        40917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        default:
        begin
            RED=8'h00;
            GRN=8'h00;
            BLU=8'h00;
        end
     endcase
endmodule