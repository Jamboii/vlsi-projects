`timescale 1ns / 1ps
module paddle_120x40_rom(
    input  [6:0] x_idx,
    input  [5:0] y_idx,
    output reg [7:0] RED,
    output reg [7:0] GRN,
    output reg [7:0] BLU);
always @ (*)
    case ({y_idx,x_idx})
        0:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        2:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        3:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        6:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        7:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        8:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        9:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        10:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        11:
        begin
            RED=8'd22;
            GRN=8'd25;
            BLU=8'd72;
        end
        12:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        13:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        14:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        15:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        16:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        17:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        18:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        19:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        20:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        21:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        22:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        23:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        24:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        25:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        26:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        27:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        28:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        29:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        30:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        31:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        32:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        33:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        34:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        35:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        36:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        37:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        38:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        39:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        40:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        41:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        42:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        43:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        44:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        45:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        46:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        47:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        48:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        49:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        50:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        51:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        52:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        53:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        54:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        55:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        56:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        57:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        58:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        59:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        60:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        61:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        62:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        63:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        64:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        65:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        66:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        67:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        68:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        69:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        70:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        71:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        72:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        73:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        74:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        75:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        76:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        77:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        78:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        79:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        80:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        81:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        82:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        83:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        84:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        85:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        86:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        87:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        88:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        89:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        90:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        91:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        92:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        93:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        94:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        95:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        96:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        97:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        98:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        99:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        100:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        101:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        102:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        103:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        104:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        105:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        106:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        107:
        begin
            RED=8'd31;
            GRN=8'd35;
            BLU=8'd99;
        end
        108:
        begin
            RED=8'd22;
            GRN=8'd25;
            BLU=8'd72;
        end
        109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        112:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        113:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        114:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        115:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        116:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        117:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        118:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        119:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        128:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        129:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        130:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        131:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        132:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        133:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        134:
        begin
            RED=8'd8;
            GRN=8'd10;
            BLU=8'd27;
        end
        135:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        136:
        begin
            RED=8'd42;
            GRN=8'd48;
            BLU=8'd137;
        end
        137:
        begin
            RED=8'd61;
            GRN=8'd70;
            BLU=8'd199;
        end
        138:
        begin
            RED=8'd61;
            GRN=8'd70;
            BLU=8'd199;
        end
        139:
        begin
            RED=8'd63;
            GRN=8'd71;
            BLU=8'd203;
        end
        140:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        141:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        142:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        143:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        144:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        145:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        146:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        147:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        148:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        149:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        150:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        151:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        152:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        153:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        154:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        155:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        156:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        157:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        158:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        159:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        160:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        161:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        162:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        163:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        164:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        165:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        166:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        167:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        168:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        169:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        170:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        171:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        172:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        173:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        174:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        175:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        176:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        177:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        178:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        179:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        180:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        181:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        182:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        183:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        184:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        185:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        186:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        187:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        188:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        189:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        190:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        191:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        192:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        193:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        194:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        195:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        196:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        197:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        198:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        199:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        200:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        201:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        202:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        203:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        204:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        205:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        206:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        207:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        208:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        209:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        210:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        211:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        212:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        213:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        214:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        215:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        216:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        217:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        218:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        219:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        220:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        221:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        222:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        223:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        224:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        225:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        226:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        227:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        228:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        229:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        230:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        231:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        232:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        233:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        234:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        235:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        236:
        begin
            RED=8'd63;
            GRN=8'd71;
            BLU=8'd203;
        end
        237:
        begin
            RED=8'd61;
            GRN=8'd70;
            BLU=8'd199;
        end
        238:
        begin
            RED=8'd61;
            GRN=8'd70;
            BLU=8'd199;
        end
        239:
        begin
            RED=8'd42;
            GRN=8'd48;
            BLU=8'd137;
        end
        240:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        241:
        begin
            RED=8'd8;
            GRN=8'd10;
            BLU=8'd27;
        end
        242:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        243:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        244:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        245:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        246:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        247:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        256:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        257:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        258:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        259:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        260:
        begin
            RED=8'd27;
            GRN=8'd31;
            BLU=8'd87;
        end
        261:
        begin
            RED=8'd48;
            GRN=8'd54;
            BLU=8'd155;
        end
        262:
        begin
            RED=8'd61;
            GRN=8'd69;
            BLU=8'd197;
        end
        263:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        264:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        265:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        266:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        267:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        268:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        269:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        270:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        271:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        272:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        273:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        274:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        275:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        276:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        277:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        278:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        279:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        280:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        281:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        282:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        283:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        284:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        285:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        286:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        287:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        288:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        289:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        290:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        291:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        292:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        293:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        294:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        295:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        296:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        297:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        298:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        299:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        300:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        301:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        302:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        303:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        304:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        305:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        306:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        307:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        308:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        309:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        310:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        311:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        312:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        313:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        314:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        315:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        316:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        317:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        318:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        319:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        320:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        321:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        322:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        323:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        324:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        325:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        326:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        327:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        328:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        329:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        330:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        331:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        332:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        333:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        334:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        335:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        336:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        337:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        338:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        339:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        340:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        341:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        342:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        343:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        344:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        345:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        346:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        347:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        348:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        349:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        350:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        351:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        352:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        353:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        354:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        355:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        356:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        357:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        358:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        359:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        360:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        361:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        362:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        363:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        364:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        365:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        366:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        367:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        368:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        369:
        begin
            RED=8'd61;
            GRN=8'd69;
            BLU=8'd197;
        end
        370:
        begin
            RED=8'd48;
            GRN=8'd54;
            BLU=8'd155;
        end
        371:
        begin
            RED=8'd27;
            GRN=8'd31;
            BLU=8'd87;
        end
        372:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        373:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        374:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        375:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        384:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        385:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        386:
        begin
            RED=8'd15;
            GRN=8'd17;
            BLU=8'd49;
        end
        387:
        begin
            RED=8'd51;
            GRN=8'd58;
            BLU=8'd165;
        end
        388:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        389:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        390:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        391:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        392:
        begin
            RED=8'd95;
            GRN=8'd101;
            BLU=8'd170;
        end
        393:
        begin
            RED=8'd142;
            GRN=8'd142;
            BLU=8'd120;
        end
        394:
        begin
            RED=8'd79;
            GRN=8'd86;
            BLU=8'd187;
        end
        395:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        396:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        397:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        398:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        399:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        400:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        401:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        402:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        403:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        404:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        405:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        406:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        407:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        408:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        409:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        410:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        411:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        412:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        413:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        414:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        415:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        416:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        417:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        418:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        419:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        420:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        421:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        422:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        423:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        424:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        425:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        426:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        427:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        428:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        429:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        430:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        431:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        432:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        433:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        434:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        435:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        436:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        437:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        438:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        439:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        440:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        441:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        442:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        443:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        444:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        445:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        446:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        447:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        448:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        449:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        450:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        451:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        452:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        453:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        454:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        455:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        456:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        457:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        458:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        459:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        460:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        461:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        462:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        463:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        464:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        465:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        466:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        467:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        468:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        469:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        470:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        471:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        472:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        473:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        474:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        475:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        476:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        477:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        478:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        479:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        480:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        481:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        482:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        483:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        484:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        485:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        486:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        487:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        488:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        489:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        490:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        491:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        492:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        493:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        494:
        begin
            RED=8'd116;
            GRN=8'd118;
            BLU=8'd148;
        end
        495:
        begin
            RED=8'd95;
            GRN=8'd101;
            BLU=8'd170;
        end
        496:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        497:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        498:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        499:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        500:
        begin
            RED=8'd58;
            GRN=8'd66;
            BLU=8'd188;
        end
        501:
        begin
            RED=8'd17;
            GRN=8'd19;
            BLU=8'd54;
        end
        502:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        503:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        512:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        513:
        begin
            RED=8'd14;
            GRN=8'd15;
            BLU=8'd43;
        end
        514:
        begin
            RED=8'd60;
            GRN=8'd69;
            BLU=8'd195;
        end
        515:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        516:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        517:
        begin
            RED=8'd110;
            GRN=8'd113;
            BLU=8'd154;
        end
        518:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        519:
        begin
            RED=8'd235;
            GRN=8'd225;
            BLU=8'd21;
        end
        520:
        begin
            RED=8'd243;
            GRN=8'd232;
            BLU=8'd12;
        end
        521:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        522:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        523:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        524:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        525:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        526:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        527:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        528:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        529:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        530:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        531:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        532:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        533:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        534:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        535:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        536:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        537:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        538:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        539:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        540:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        541:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        542:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        543:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        544:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        545:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        546:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        547:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        548:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        549:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        550:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        551:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        552:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        553:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        554:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        555:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        556:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        557:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        558:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        559:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        560:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        561:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        562:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        563:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        564:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        565:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        566:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        567:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        568:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        569:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        570:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        571:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        572:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        573:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        574:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        575:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        576:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        577:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        578:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        579:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        580:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        581:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        582:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        583:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        584:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        585:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        586:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        587:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        588:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        589:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        590:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        591:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        592:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        593:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        594:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        595:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        596:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        597:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        598:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        599:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        600:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        601:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        602:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        603:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        604:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        605:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        606:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        607:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        608:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        609:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        610:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        611:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        612:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        613:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        614:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        615:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        616:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        617:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        618:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        619:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        620:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        621:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        622:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        623:
        begin
            RED=8'd243;
            GRN=8'd232;
            BLU=8'd12;
        end
        624:
        begin
            RED=8'd235;
            GRN=8'd225;
            BLU=8'd21;
        end
        625:
        begin
            RED=8'd165;
            GRN=8'd163;
            BLU=8'd95;
        end
        626:
        begin
            RED=8'd110;
            GRN=8'd113;
            BLU=8'd154;
        end
        627:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        628:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        629:
        begin
            RED=8'd60;
            GRN=8'd69;
            BLU=8'd195;
        end
        630:
        begin
            RED=8'd20;
            GRN=8'd23;
            BLU=8'd64;
        end
        631:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        640:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        641:
        begin
            RED=8'd54;
            GRN=8'd62;
            BLU=8'd175;
        end
        642:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        643:
        begin
            RED=8'd98;
            GRN=8'd103;
            BLU=8'd167;
        end
        644:
        begin
            RED=8'd201;
            GRN=8'd195;
            BLU=8'd57;
        end
        645:
        begin
            RED=8'd246;
            GRN=8'd234;
            BLU=8'd10;
        end
        646:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        647:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        648:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        649:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        650:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        651:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        652:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        653:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        654:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        655:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        656:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        657:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        658:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        659:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        660:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        661:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        662:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        663:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        664:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        665:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        666:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        667:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        668:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        669:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        670:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        671:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        672:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        673:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        674:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        675:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        676:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        677:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        678:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        679:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        680:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        681:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        682:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        683:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        684:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        685:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        686:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        687:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        688:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        689:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        690:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        691:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        692:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        693:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        694:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        695:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        696:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        697:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        698:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        699:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        700:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        701:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        702:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        703:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        704:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        705:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        706:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        707:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        708:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        709:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        710:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        711:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        712:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        713:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        714:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        715:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        716:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        717:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        718:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        719:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        720:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        721:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        722:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        723:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        724:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        725:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        726:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        727:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        728:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        729:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        730:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        731:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        732:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        733:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        734:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        735:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        736:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        737:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        738:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        739:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        740:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        741:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        742:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        743:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        744:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        745:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        746:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        747:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        748:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        749:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        750:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        751:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        752:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        753:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        754:
        begin
            RED=8'd246;
            GRN=8'd234;
            BLU=8'd10;
        end
        755:
        begin
            RED=8'd201;
            GRN=8'd195;
            BLU=8'd57;
        end
        756:
        begin
            RED=8'd116;
            GRN=8'd119;
            BLU=8'd147;
        end
        757:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        758:
        begin
            RED=8'd58;
            GRN=8'd66;
            BLU=8'd187;
        end
        759:
        begin
            RED=8'd4;
            GRN=8'd5;
            BLU=8'd14;
        end
        768:
        begin
            RED=8'd10;
            GRN=8'd12;
            BLU=8'd34;
        end
        769:
        begin
            RED=8'd62;
            GRN=8'd71;
            BLU=8'd202;
        end
        770:
        begin
            RED=8'd132;
            GRN=8'd133;
            BLU=8'd132;
        end
        771:
        begin
            RED=8'd241;
            GRN=8'd229;
            BLU=8'd15;
        end
        772:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        773:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        774:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        775:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        776:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        777:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        778:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        779:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        780:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        781:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        782:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        783:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        784:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        785:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        786:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        787:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        788:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        789:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        790:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        791:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        792:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        793:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        794:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        795:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        796:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        797:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        798:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        799:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        800:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        801:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        802:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        803:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        804:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        805:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        806:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        807:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        808:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        809:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        810:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        811:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        812:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        813:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        814:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        815:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        816:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        817:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        818:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        819:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        820:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        821:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        822:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        823:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        824:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        825:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        826:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        827:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        828:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        829:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        830:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        831:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        832:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        833:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        834:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        835:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        836:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        837:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        838:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        839:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        840:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        841:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        842:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        843:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        844:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        845:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        846:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        847:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        848:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        849:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        850:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        851:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        852:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        853:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        854:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        855:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        856:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        857:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        858:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        859:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        860:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        861:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        862:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        863:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        864:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        865:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        866:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        867:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        868:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        869:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        870:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        871:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        872:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        873:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        874:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        875:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        876:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        877:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        878:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        879:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        880:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        881:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        882:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        883:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        884:
        begin
            RED=8'd248;
            GRN=8'd236;
            BLU=8'd7;
        end
        885:
        begin
            RED=8'd149;
            GRN=8'd148;
            BLU=8'd113;
        end
        886:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        887:
        begin
            RED=8'd18;
            GRN=8'd20;
            BLU=8'd58;
        end
        896:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        897:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        898:
        begin
            RED=8'd218;
            GRN=8'd209;
            BLU=8'd40;
        end
        899:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        900:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        901:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        902:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        903:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        904:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        905:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        906:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        907:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        908:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        909:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        910:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        911:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        912:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        913:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        914:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        915:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        916:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        917:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        918:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        919:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        920:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        921:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        922:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        923:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        924:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        925:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        926:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        927:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        928:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        929:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        930:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        931:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        932:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        933:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        934:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        935:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        936:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        937:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        938:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        939:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        940:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        941:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        942:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        943:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        944:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        945:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        946:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        947:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        948:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        949:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        950:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        951:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        952:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        953:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        954:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        955:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        956:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        957:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        958:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        959:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        960:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        961:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        962:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        963:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        964:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        965:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        966:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        967:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        968:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        969:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        970:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        971:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        972:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        973:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        974:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        975:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        976:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        977:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        978:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        979:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        980:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        981:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        982:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        983:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        984:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        985:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        986:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        987:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        988:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        989:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        990:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        991:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        992:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        993:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        994:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        995:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        996:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        997:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        998:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        999:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1000:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1001:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1002:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1003:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1004:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1005:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1006:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        1007:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1008:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1009:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1010:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1011:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1012:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1013:
        begin
            RED=8'd250;
            GRN=8'd238;
            BLU=8'd5;
        end
        1014:
        begin
            RED=8'd82;
            GRN=8'd89;
            BLU=8'd183;
        end
        1015:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        1024:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        1025:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1026:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        1027:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1028:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1029:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1030:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1031:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1032:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1033:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1034:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        1035:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1036:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1037:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1038:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1039:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1040:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1041:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1042:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1043:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1044:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1045:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1046:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1047:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1048:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1049:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1050:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1051:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1052:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1053:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1054:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1055:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1056:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1057:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1058:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1059:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1060:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1061:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1062:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1063:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1064:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1065:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1066:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1067:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1068:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1069:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1070:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1071:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1072:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1073:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1074:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1075:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1076:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1077:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1078:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1079:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1080:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1081:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1082:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1083:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1084:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1085:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1086:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1087:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1088:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1089:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1090:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1091:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1092:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1093:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1094:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1095:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1096:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1097:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1098:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1099:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1100:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1101:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1102:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1103:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1104:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1105:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1106:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1107:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1108:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1109:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1110:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1111:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1112:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1113:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1114:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1115:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1116:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1117:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1118:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1119:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1120:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1121:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1122:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1123:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1124:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1125:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1126:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1127:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1128:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1129:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1130:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1131:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1132:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1133:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1134:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        1135:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1136:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1137:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1138:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1139:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1140:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1141:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1142:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        1143:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        1152:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        1153:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1154:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        1155:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1156:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1157:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1158:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1159:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1160:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1161:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1162:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        1163:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1164:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1165:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1166:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1167:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1168:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1169:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1170:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1171:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1172:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1173:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1174:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1175:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1176:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1177:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1178:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1179:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1180:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1181:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1182:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1183:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1184:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1185:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1186:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1187:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1188:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1189:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1190:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1191:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1192:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1193:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1194:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1195:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1196:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1197:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1198:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1199:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1200:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1201:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1202:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1203:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1204:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1205:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1206:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1207:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1208:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1209:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1210:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1211:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1212:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1213:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1214:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1215:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1216:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1217:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1218:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1219:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1220:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1221:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1222:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1223:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1224:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1225:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1226:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1227:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1228:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1229:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1230:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1231:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1232:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1233:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1234:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1235:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1236:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1237:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1238:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1239:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1240:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1241:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1242:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1243:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1244:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1245:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1246:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1247:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1248:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1249:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1250:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1251:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1252:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1253:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1254:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1255:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1256:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1257:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1258:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1259:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1260:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1261:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1262:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        1263:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1264:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1265:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1266:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1267:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1268:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1269:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1270:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        1271:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        1280:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        1281:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1282:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        1283:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1284:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1285:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1286:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1287:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1288:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1289:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1290:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        1291:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1292:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1293:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1294:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1295:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1296:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1297:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1298:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1299:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1300:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1301:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1302:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1303:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1304:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1305:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1306:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1307:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1308:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1309:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1310:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1311:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1312:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1313:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1314:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1315:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1316:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1317:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1318:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1319:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1320:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1321:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1322:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1323:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1324:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1325:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1326:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1327:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1328:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1329:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1330:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1331:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1332:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1333:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1334:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1335:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1336:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1337:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1338:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1339:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1340:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1341:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1342:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1343:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1344:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1345:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1346:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1347:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1348:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1349:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1350:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1351:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1352:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1353:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1354:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1355:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1356:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1357:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1358:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1359:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1360:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1361:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1362:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1363:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1364:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1365:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1366:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1367:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1368:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1369:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1370:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1371:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1372:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1373:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1374:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1375:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1376:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1377:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1378:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1379:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1380:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1381:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1382:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1383:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1384:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1385:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1386:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1387:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1388:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1389:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1390:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        1391:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1392:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1393:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1394:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1395:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1396:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1397:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1398:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        1399:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        1408:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        1409:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1410:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        1411:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1412:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1413:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1414:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1415:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1416:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1417:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1418:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        1419:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1420:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1421:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1422:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1423:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1424:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1425:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1426:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1427:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1428:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1429:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1430:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1431:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1432:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1433:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1434:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1435:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1436:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1437:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1438:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1439:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1440:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1441:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1442:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1443:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1444:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1445:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1446:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1447:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1448:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1449:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1450:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1451:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1452:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1453:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1454:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1455:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1456:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1457:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1458:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1459:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1460:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1461:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1462:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1463:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1464:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1465:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1466:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1467:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1468:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1469:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1470:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1471:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1472:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1473:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1474:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1475:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1476:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1477:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1478:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1479:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1480:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1481:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1482:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1483:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1484:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1485:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1486:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1487:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1488:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1489:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1490:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1491:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1492:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1493:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1494:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1495:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1496:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1497:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1498:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1499:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1500:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1501:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1502:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1503:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1504:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1505:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1506:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1507:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1508:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1509:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1510:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1511:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1512:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1513:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1514:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1515:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1516:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1517:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1518:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        1519:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1520:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1521:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1522:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1523:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1524:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1525:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1526:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        1527:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        1536:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        1537:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1538:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        1539:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1540:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1541:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1542:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1543:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1544:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1545:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1546:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        1547:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1548:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1549:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1550:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1551:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1552:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1553:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1554:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1555:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1556:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1557:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1558:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1559:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1560:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1561:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1562:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1563:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1564:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1565:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1566:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1567:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1568:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1569:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1570:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1571:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1572:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1573:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1574:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1575:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1576:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1577:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1578:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1579:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1580:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1581:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1582:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1583:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1584:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1585:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1586:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1587:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1588:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1589:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1590:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1591:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1592:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1593:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1594:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1595:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1596:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1597:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1598:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1599:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1600:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1601:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1602:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1603:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1604:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1605:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1606:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1607:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1608:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1609:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1610:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1611:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1612:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1613:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1614:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1615:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1616:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1617:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1618:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1619:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1620:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1621:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1622:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1623:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1624:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1625:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1626:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1627:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1628:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1629:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1630:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1631:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1632:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1633:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1634:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1635:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1636:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1637:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1638:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1639:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1640:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1641:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1642:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1643:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1644:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1645:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1646:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        1647:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1648:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1649:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1650:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1651:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1652:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1653:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1654:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        1655:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        1664:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        1665:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1666:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        1667:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1668:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1669:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1670:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1671:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1672:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1673:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1674:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        1675:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1676:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1677:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1678:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1679:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1680:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1681:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1682:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1683:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1684:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1685:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1686:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1687:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1688:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1689:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1690:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1691:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1692:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1693:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1694:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1695:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1696:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1697:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1698:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1699:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1700:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1701:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1702:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1703:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1704:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1705:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1706:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1707:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1708:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1709:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1710:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1711:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1712:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1713:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1714:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1715:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1716:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1717:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1718:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1719:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1720:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1721:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1722:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1723:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1724:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1725:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1726:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1727:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1728:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1729:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1730:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1731:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1732:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1733:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1734:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1735:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1736:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1737:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1738:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1739:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1740:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1741:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1742:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1743:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1744:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1745:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1746:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1747:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1748:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1749:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1750:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1751:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1752:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1753:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1754:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1755:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1756:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1757:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1758:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1759:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1760:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1761:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1762:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1763:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1764:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1765:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1766:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1767:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1768:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1769:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1770:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1771:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1772:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1773:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1774:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        1775:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1776:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1777:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1778:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1779:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1780:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1781:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1782:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        1783:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        1792:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        1793:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1794:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        1795:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1796:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1797:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1798:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1799:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1800:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1801:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1802:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        1803:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1804:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1805:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1806:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1807:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1808:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1809:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1810:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1811:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1812:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1813:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1814:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1815:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1816:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1817:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1818:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1819:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1820:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1821:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1822:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1823:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1824:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1825:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1826:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1827:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1828:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1829:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1830:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1831:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1832:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1833:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1834:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1835:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1836:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1837:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1838:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1839:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1840:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1841:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1842:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1843:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1844:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1845:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1846:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1847:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1848:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1849:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1850:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1851:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1852:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1853:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1854:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1855:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1856:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1857:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1858:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1859:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1860:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1861:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1862:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1863:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1864:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1865:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1866:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1867:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1868:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1869:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1870:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1871:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1872:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1873:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1874:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1875:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1876:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1877:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1878:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1879:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1880:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1881:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1882:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1883:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1884:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1885:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1886:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1887:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1888:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1889:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1890:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1891:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1892:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1893:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1894:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1895:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1896:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1897:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1898:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1899:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1900:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1901:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1902:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        1903:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1904:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1905:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1906:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1907:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1908:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1909:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1910:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        1911:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        1920:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        1921:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1922:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        1923:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1924:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1925:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1926:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1927:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1928:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1929:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        1930:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        1931:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1932:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1933:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1934:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1935:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1936:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1937:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1938:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1939:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1940:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1941:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1942:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1943:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1944:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1945:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1946:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1947:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1948:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1949:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1950:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1951:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1952:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1953:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1954:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1955:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1956:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1957:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1958:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1959:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1960:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1961:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1962:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1963:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1964:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1965:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1966:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1967:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1968:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1969:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1970:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1971:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1972:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1973:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1974:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1975:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1976:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1977:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1978:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1979:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1980:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1981:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1982:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1983:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1984:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1985:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1986:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1987:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1988:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1989:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1990:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1991:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1992:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1993:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1994:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1995:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1996:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1997:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1998:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        1999:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2000:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2001:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2002:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2003:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2004:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2005:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2006:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2007:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2008:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2009:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2010:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2011:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2012:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2013:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2014:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2015:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2016:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2017:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2018:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2019:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2020:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2021:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2022:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2023:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2024:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2025:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2026:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2027:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2028:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2029:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2030:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        2031:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2032:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2033:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2034:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2035:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2036:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2037:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2038:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        2039:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        2048:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        2049:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2050:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        2051:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2052:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2053:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2054:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2055:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2056:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2057:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2058:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        2059:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2060:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2061:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2062:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2063:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2064:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2065:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2066:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2067:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2068:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2069:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2070:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2071:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2072:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2073:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2074:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2075:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2076:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2077:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2078:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2079:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2080:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2081:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2082:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2083:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2084:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2085:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2086:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2087:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2088:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2089:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2090:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2091:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2092:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2093:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2094:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2095:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2096:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2097:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2098:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2099:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2100:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2101:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2102:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2103:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2104:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2105:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2106:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2107:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2108:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2109:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2110:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2111:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2112:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2113:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2114:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2115:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2116:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2117:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2118:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2119:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2120:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2121:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2122:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2123:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2124:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2125:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2126:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2127:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2128:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2129:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2130:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2131:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2132:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2133:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2134:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2135:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2136:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2137:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2138:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2139:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2140:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2141:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2142:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2143:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2144:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2145:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2146:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2147:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2148:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2149:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2150:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2151:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2152:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2153:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2154:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2155:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2156:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2157:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2158:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        2159:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2160:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2161:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2162:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2163:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2164:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2165:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2166:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        2167:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        2176:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        2177:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2178:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        2179:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2180:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2181:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2182:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2183:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2184:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2185:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2186:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        2187:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2188:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2189:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2190:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2191:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2192:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2193:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2194:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2195:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2196:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2197:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2198:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2199:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2200:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2201:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2202:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2203:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2204:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2205:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2206:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2207:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2208:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2209:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2210:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2211:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2212:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2213:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2214:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2215:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2216:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2217:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2218:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2219:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2220:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2221:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2222:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2223:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2224:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2225:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2226:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2227:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2228:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2229:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2230:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2231:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2232:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2233:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2234:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2235:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2236:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2237:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2238:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2239:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2240:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2241:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2242:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2243:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2244:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2245:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2246:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2247:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2248:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2249:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2250:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2251:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2252:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2253:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2254:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2255:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2256:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2257:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2258:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2259:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2260:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2261:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2262:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2263:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2264:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2265:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2266:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2267:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2268:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2269:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2270:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2271:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2272:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2273:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2274:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2275:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2276:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2277:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2278:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2279:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2280:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2281:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2282:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2283:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2284:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2285:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2286:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        2287:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2288:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2289:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2290:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2291:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2292:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2293:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2294:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        2295:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        2304:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        2305:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2306:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        2307:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2308:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2309:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2310:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2311:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2312:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2313:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2314:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        2315:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2316:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2317:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2318:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2319:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2320:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2321:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2322:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2323:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2324:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2325:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2326:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2327:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2328:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2329:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2330:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2331:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2332:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2333:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2334:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2335:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2336:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2337:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2338:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2339:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2340:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2341:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2342:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2343:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2344:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2345:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2346:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2347:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2348:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2349:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2350:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2351:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2352:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2353:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2354:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2355:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2356:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2357:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2358:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2359:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2360:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2361:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2362:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2363:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2364:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2365:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2366:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2367:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2368:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2369:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2370:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2371:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2372:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2373:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2374:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2375:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2376:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2377:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2378:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2379:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2380:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2381:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2382:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2383:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2384:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2385:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2386:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2387:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2388:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2389:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2390:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2391:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2392:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2393:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2394:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2395:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2396:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2397:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2398:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2399:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2400:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2401:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2402:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2403:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2404:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2405:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2406:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2407:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2408:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2409:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2410:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2411:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2412:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2413:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2414:
        begin
            RED=8'd191;
            GRN=8'd185;
            BLU=8'd68;
        end
        2415:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2416:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2417:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2418:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2419:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2420:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2421:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2422:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        2423:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        2432:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        2433:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2434:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        2435:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2436:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2437:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2438:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2439:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2440:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2441:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2442:
        begin
            RED=8'd102;
            GRN=8'd106;
            BLU=8'd163;
        end
        2443:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2444:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2445:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2446:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2447:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2448:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2449:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2450:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2451:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2452:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2453:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2454:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2455:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2456:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2457:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2458:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2459:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2460:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2461:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2462:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2463:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2464:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2465:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2466:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2467:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2468:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2469:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2470:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2471:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2472:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2473:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2474:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2475:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2476:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2477:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2478:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2479:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2480:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2481:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2482:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2483:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2484:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2485:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2486:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2487:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2488:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2489:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2490:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2491:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2492:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2493:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2494:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2495:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2496:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2497:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2498:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2499:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2500:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2501:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2502:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2503:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2504:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2505:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2506:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2507:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2508:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2509:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2510:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2511:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2512:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2513:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2514:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2515:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2516:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2517:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2518:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2519:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2520:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2521:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2522:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2523:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2524:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2525:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2526:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2527:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2528:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2529:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2530:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2531:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2532:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2533:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2534:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2535:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2536:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2537:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2538:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2539:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2540:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2541:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2542:
        begin
            RED=8'd164;
            GRN=8'd161;
            BLU=8'd96;
        end
        2543:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2544:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2545:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2546:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2547:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2548:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2549:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2550:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        2551:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        2560:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        2561:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2562:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        2563:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2564:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2565:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2566:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2567:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2568:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2569:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2570:
        begin
            RED=8'd127;
            GRN=8'd128;
            BLU=8'd136;
        end
        2571:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2572:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2573:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2574:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2575:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2576:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2577:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2578:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2579:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2580:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2581:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2582:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2583:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2584:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2585:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2586:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2587:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2588:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2589:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2590:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2591:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2592:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2593:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2594:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2595:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2596:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2597:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2598:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2599:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2600:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2601:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2602:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2603:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2604:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2605:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2606:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2607:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2608:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2609:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2610:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2611:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2612:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2613:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2614:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2615:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2616:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2617:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2618:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2619:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2620:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2621:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2622:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2623:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2624:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2625:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2626:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2627:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2628:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2629:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2630:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2631:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2632:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2633:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2634:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2635:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2636:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2637:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2638:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2639:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2640:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2641:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2642:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2643:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2644:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2645:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2646:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2647:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2648:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2649:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2650:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2651:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2652:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2653:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2654:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2655:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2656:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2657:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2658:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2659:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2660:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2661:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2662:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2663:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2664:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2665:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2666:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2667:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2668:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2669:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2670:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        2671:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2672:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2673:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2674:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2675:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2676:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2677:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2678:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        2679:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        2688:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        2689:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2690:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        2691:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2692:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2693:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2694:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2695:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2696:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2697:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2698:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        2699:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2700:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2701:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2702:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2703:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2704:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2705:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2706:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2707:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2708:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2709:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2710:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2711:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2712:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2713:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2714:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2715:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2716:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2717:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2718:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2719:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2720:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2721:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2722:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2723:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2724:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2725:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2726:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2727:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2728:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2729:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2730:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2731:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2732:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2733:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2734:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2735:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2736:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2737:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2738:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2739:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2740:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2741:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2742:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2743:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2744:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2745:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2746:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2747:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2748:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2749:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2750:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2751:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2752:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2753:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2754:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2755:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2756:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2757:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2758:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2759:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2760:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2761:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2762:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2763:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2764:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2765:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2766:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2767:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2768:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2769:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2770:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2771:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2772:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2773:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2774:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2775:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2776:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2777:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2778:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2779:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2780:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2781:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2782:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2783:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2784:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2785:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2786:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2787:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2788:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2789:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2790:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2791:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2792:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2793:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2794:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2795:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2796:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2797:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2798:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        2799:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2800:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2801:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2802:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2803:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2804:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2805:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2806:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        2807:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        2816:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        2817:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2818:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        2819:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2820:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2821:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2822:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2823:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2824:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2825:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2826:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        2827:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2828:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2829:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2830:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2831:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2832:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2833:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2834:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2835:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2836:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2837:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2838:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2839:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2840:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2841:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2842:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2843:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2844:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2845:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2846:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2847:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2848:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2849:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2850:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2851:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2852:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2853:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2854:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2855:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2856:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2857:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2858:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2859:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2860:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2861:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2862:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2863:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2864:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2865:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2866:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2867:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2868:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2869:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2870:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2871:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2872:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2873:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2874:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2875:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2876:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2877:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2878:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2879:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2880:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2881:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2882:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2883:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2884:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2885:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2886:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2887:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2888:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2889:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2890:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2891:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2892:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2893:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2894:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2895:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2896:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2897:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2898:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2899:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2900:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2901:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2902:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2903:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2904:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2905:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2906:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2907:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2908:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2909:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2910:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2911:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2912:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2913:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2914:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2915:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2916:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2917:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2918:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2919:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2920:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2921:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2922:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2923:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2924:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2925:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2926:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        2927:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2928:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2929:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2930:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2931:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2932:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2933:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2934:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        2935:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        2944:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        2945:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2946:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        2947:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2948:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2949:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2950:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2951:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2952:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2953:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        2954:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        2955:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2956:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2957:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2958:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2959:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2960:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2961:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2962:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2963:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2964:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2965:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2966:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2967:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2968:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2969:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2970:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2971:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2972:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2973:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2974:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2975:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2976:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2977:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2978:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2979:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2980:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2981:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2982:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2983:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2984:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2985:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2986:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2987:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2988:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2989:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2990:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2991:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2992:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2993:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2994:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2995:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2996:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2997:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2998:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        2999:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3000:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3001:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3002:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3003:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3004:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3005:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3006:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3007:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3008:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3009:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3010:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3011:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3012:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3013:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3014:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3015:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3016:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3017:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3018:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3019:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3020:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3021:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3022:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3023:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3024:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3025:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3026:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3027:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3028:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3029:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3030:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3031:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3032:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3033:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3034:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3035:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3036:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3037:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3038:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3039:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3040:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3041:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3042:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3043:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3044:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3045:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3046:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3047:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3048:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3049:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3050:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3051:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3052:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3053:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3054:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        3055:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3056:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3057:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3058:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3059:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3060:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3061:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3062:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        3063:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        3072:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        3073:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3074:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        3075:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3076:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3077:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3078:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3079:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3080:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3081:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3082:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        3083:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3084:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3085:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3086:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3087:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3088:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3089:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3090:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3091:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3092:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3093:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3094:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3095:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3096:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3097:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3098:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3099:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3100:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3101:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3102:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3103:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3104:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3105:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3106:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3107:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3108:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3109:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3110:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3111:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3112:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3113:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3114:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3115:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3116:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3117:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3118:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3119:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3120:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3121:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3122:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3123:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3124:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3125:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3126:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3127:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3128:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3129:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3130:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3131:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3132:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3133:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3134:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3135:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3136:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3137:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3138:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3139:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3140:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3141:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3142:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3143:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3144:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3145:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3146:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3147:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3148:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3149:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3150:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3151:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3152:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3153:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3154:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3155:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3156:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3157:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3158:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3159:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3160:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3161:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3162:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3163:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3164:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3165:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3166:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3167:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3168:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3169:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3170:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3171:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3172:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3173:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3174:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3175:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3176:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3177:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3178:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3179:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3180:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3181:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3182:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        3183:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3184:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3185:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3186:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3187:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3188:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3189:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3190:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        3191:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        3200:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        3201:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3202:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        3203:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3204:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3205:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3206:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3207:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3208:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3209:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3210:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        3211:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3212:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3213:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3214:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3215:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3216:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3217:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3218:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3219:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3220:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3221:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3222:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3223:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3224:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3225:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3226:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3227:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3228:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3229:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3230:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3231:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3232:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3233:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3234:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3235:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3236:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3237:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3238:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3239:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3240:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3241:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3242:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3243:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3244:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3245:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3246:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3247:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3248:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3249:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3250:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3251:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3252:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3253:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3254:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3255:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3256:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3257:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3258:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3259:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3260:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3261:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3262:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3263:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3264:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3265:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3266:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3267:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3268:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3269:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3270:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3271:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3272:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3273:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3274:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3275:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3276:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3277:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3278:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3279:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3280:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3281:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3282:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3283:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3284:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3285:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3286:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3287:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3288:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3289:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3290:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3291:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3292:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3293:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3294:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3295:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3296:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3297:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3298:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3299:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3300:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3301:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3302:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3303:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3304:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3305:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3306:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3307:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3308:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3309:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3310:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        3311:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3312:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3313:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3314:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3315:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3316:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3317:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3318:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        3319:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        3328:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        3329:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3330:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        3331:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3332:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3333:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3334:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3335:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3336:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3337:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3338:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        3339:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3340:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3341:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3342:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3343:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3344:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3345:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3346:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3347:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3348:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3349:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3350:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3351:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3352:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3353:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3354:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3355:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3356:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3357:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3358:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3359:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3360:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3361:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3362:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3363:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3364:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3365:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3366:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3367:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3368:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3369:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3370:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3371:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3372:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3373:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3374:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3375:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3376:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3377:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3378:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3379:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3380:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3381:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3382:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3383:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3384:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3385:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3386:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3387:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3388:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3389:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3390:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3391:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3392:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3393:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3394:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3395:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3396:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3397:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3398:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3399:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3400:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3401:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3402:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3403:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3404:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3405:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3406:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3407:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3408:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3409:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3410:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3411:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3412:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3413:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3414:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3415:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3416:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3417:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3418:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3419:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3420:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3421:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3422:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3423:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3424:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3425:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3426:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3427:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3428:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3429:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3430:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3431:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3432:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3433:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3434:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3435:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3436:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3437:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3438:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        3439:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3440:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3441:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3442:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3443:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3444:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3445:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3446:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        3447:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        3456:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        3457:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3458:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        3459:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3460:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3461:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3462:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3463:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3464:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3465:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3466:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        3467:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3468:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3469:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3470:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3471:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3472:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3473:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3474:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3475:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3476:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3477:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3478:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3479:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3480:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3481:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3482:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3483:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3484:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3485:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3486:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3487:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3488:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3489:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3490:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3491:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3492:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3493:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3494:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3495:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3496:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3497:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3498:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3499:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3500:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3501:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3502:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3503:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3504:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3505:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3506:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3507:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3508:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3509:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3510:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3511:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3512:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3513:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3514:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3515:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3516:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3517:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3518:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3519:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3520:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3521:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3522:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3523:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3524:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3525:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3526:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3527:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3528:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3529:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3530:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3531:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3532:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3533:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3534:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3535:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3536:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3537:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3538:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3539:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3540:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3541:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3542:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3543:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3544:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3545:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3546:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3547:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3548:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3549:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3550:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3551:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3552:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3553:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3554:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3555:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3556:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3557:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3558:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3559:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3560:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3561:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3562:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3563:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3564:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3565:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3566:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        3567:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3568:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3569:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3570:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3571:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3572:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3573:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3574:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        3575:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        3584:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        3585:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3586:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        3587:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3588:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3589:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3590:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3591:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3592:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3593:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3594:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        3595:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3596:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3597:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3598:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3599:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3600:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3601:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3602:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3603:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3604:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3605:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3606:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3607:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3608:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3609:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3610:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3611:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3612:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3613:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3614:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3615:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3616:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3617:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3618:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3619:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3620:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3621:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3622:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3623:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3624:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3625:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3626:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3627:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3628:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3629:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3630:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3631:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3632:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3633:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3634:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3635:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3636:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3637:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3638:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3639:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3640:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3641:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3642:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3643:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3644:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3645:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3646:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3647:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3648:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3649:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3650:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3651:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3652:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3653:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3654:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3655:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3656:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3657:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3658:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3659:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3660:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3661:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3662:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3663:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3664:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3665:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3666:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3667:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3668:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3669:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3670:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3671:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3672:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3673:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3674:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3675:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3676:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3677:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3678:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3679:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3680:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3681:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3682:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3683:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3684:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3685:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3686:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3687:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3688:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3689:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3690:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3691:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3692:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3693:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3694:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        3695:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3696:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3697:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3698:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3699:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3700:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3701:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3702:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        3703:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        3712:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        3713:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3714:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        3715:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3716:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3717:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3718:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3719:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3720:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3721:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3722:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        3723:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3724:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3725:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3726:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3727:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3728:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3729:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3730:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3731:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3732:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3733:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3734:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3735:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3736:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3737:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3738:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3739:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3740:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3741:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3742:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3743:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3744:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3745:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3746:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3747:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3748:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3749:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3750:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3751:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3752:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3753:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3754:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3755:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3756:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3757:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3758:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3759:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3760:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3761:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3762:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3763:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3764:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3765:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3766:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3767:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3768:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3769:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3770:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3771:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3772:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3773:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3774:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3775:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3776:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3777:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3778:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3779:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3780:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3781:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3782:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3783:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3784:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3785:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3786:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3787:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3788:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3789:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3790:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3791:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3792:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3793:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3794:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3795:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3796:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3797:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3798:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3799:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3800:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3801:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3802:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3803:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3804:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3805:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3806:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3807:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3808:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3809:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3810:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3811:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3812:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3813:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3814:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3815:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3816:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3817:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3818:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3819:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3820:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3821:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3822:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        3823:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3824:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3825:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3826:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3827:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3828:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3829:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3830:
        begin
            RED=8'd86;
            GRN=8'd93;
            BLU=8'd179;
        end
        3831:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        3840:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        3841:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3842:
        begin
            RED=8'd227;
            GRN=8'd217;
            BLU=8'd30;
        end
        3843:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3844:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3845:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3846:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3847:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3848:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3849:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3850:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        3851:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3852:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3853:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3854:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3855:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3856:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3857:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3858:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3859:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3860:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3861:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3862:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3863:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3864:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3865:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3866:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3867:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3868:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3869:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3870:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3871:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3872:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3873:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3874:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3875:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3876:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3877:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3878:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3879:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3880:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3881:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3882:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3883:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3884:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3885:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3886:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3887:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3888:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3889:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3890:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3891:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3892:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3893:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3894:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3895:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3896:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3897:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3898:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3899:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3900:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3901:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3902:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3903:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3904:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3905:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3906:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3907:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3908:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3909:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3910:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3911:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3912:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3913:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3914:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3915:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3916:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3917:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3918:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3919:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3920:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3921:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3922:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3923:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3924:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3925:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3926:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3927:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3928:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3929:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3930:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3931:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3932:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3933:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3934:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3935:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3936:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3937:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3938:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3939:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3940:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3941:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3942:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3943:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3944:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3945:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3946:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3947:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3948:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3949:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3950:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        3951:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3952:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3953:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3954:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3955:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3956:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3957:
        begin
            RED=8'd249;
            GRN=8'd236;
            BLU=8'd7;
        end
        3958:
        begin
            RED=8'd81;
            GRN=8'd88;
            BLU=8'd185;
        end
        3959:
        begin
            RED=8'd29;
            GRN=8'd33;
            BLU=8'd94;
        end
        3968:
        begin
            RED=8'd10;
            GRN=8'd11;
            BLU=8'd32;
        end
        3969:
        begin
            RED=8'd62;
            GRN=8'd71;
            BLU=8'd201;
        end
        3970:
        begin
            RED=8'd167;
            GRN=8'd164;
            BLU=8'd94;
        end
        3971:
        begin
            RED=8'd246;
            GRN=8'd234;
            BLU=8'd9;
        end
        3972:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3973:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3974:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3975:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3976:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3977:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        3978:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        3979:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3980:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3981:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3982:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3983:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3984:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3985:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3986:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3987:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3988:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3989:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3990:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3991:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3992:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3993:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3994:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3995:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3996:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3997:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3998:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        3999:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4000:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4001:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4002:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4003:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4004:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4005:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4006:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4007:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4008:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4009:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4010:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4011:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4012:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4013:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4014:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4015:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4016:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4017:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4018:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4019:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4020:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4021:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4022:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4023:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4024:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4025:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4026:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4027:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4028:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4029:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4030:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4031:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4032:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4033:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4034:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4035:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4036:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4037:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4038:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4039:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4040:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4041:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4042:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4043:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4044:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4045:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4046:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4047:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4048:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4049:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4050:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4051:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4052:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4053:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4054:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4055:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4056:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4057:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4058:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4059:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4060:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4061:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4062:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4063:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4064:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4065:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4066:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4067:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4068:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4069:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4070:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4071:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4072:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4073:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4074:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4075:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4076:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4077:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4078:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        4079:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4080:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4081:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4082:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4083:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4084:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4085:
        begin
            RED=8'd169;
            GRN=8'd165;
            BLU=8'd92;
        end
        4086:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4087:
        begin
            RED=8'd17;
            GRN=8'd19;
            BLU=8'd55;
        end
        4096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4097:
        begin
            RED=8'd55;
            GRN=8'd63;
            BLU=8'd179;
        end
        4098:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4099:
        begin
            RED=8'd132;
            GRN=8'd134;
            BLU=8'd130;
        end
        4100:
        begin
            RED=8'd226;
            GRN=8'd217;
            BLU=8'd31;
        end
        4101:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4102:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4103:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4104:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4105:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4106:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        4107:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4108:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4109:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4110:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4111:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4112:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4113:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4114:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4115:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4116:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4117:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4118:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4119:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4120:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4121:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4122:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4123:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4124:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4125:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4126:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4127:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4128:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4129:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4130:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4131:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4132:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4133:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4134:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4135:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4136:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4137:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4138:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4139:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4140:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4141:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4142:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4143:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4144:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4145:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4146:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4147:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4148:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4149:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4150:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4151:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4152:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4153:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4154:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4155:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4156:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4157:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4158:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4159:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4160:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4161:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4162:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4163:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4164:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4165:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4166:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4167:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4168:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4169:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4170:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4171:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4172:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4173:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4174:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4175:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4176:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4177:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4178:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4179:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4180:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4181:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4182:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4183:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4184:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4185:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4186:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4187:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4188:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4189:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4190:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4191:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4192:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4193:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4194:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4195:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4196:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4197:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4198:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4199:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4200:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4201:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4202:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4203:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4204:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4205:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4206:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        4207:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4208:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4209:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4210:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4211:
        begin
            RED=8'd226;
            GRN=8'd217;
            BLU=8'd31;
        end
        4212:
        begin
            RED=8'd146;
            GRN=8'd145;
            BLU=8'd116;
        end
        4213:
        begin
            RED=8'd66;
            GRN=8'd74;
            BLU=8'd201;
        end
        4214:
        begin
            RED=8'd62;
            GRN=8'd71;
            BLU=8'd201;
        end
        4215:
        begin
            RED=8'd10;
            GRN=8'd11;
            BLU=8'd33;
        end
        4224:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4225:
        begin
            RED=8'd26;
            GRN=8'd30;
            BLU=8'd85;
        end
        4226:
        begin
            RED=8'd62;
            GRN=8'd70;
            BLU=8'd199;
        end
        4227:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4228:
        begin
            RED=8'd74;
            GRN=8'd82;
            BLU=8'd193;
        end
        4229:
        begin
            RED=8'd127;
            GRN=8'd129;
            BLU=8'd136;
        end
        4230:
        begin
            RED=8'd208;
            GRN=8'd200;
            BLU=8'd50;
        end
        4231:
        begin
            RED=8'd232;
            GRN=8'd222;
            BLU=8'd25;
        end
        4232:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4233:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4234:
        begin
            RED=8'd153;
            GRN=8'd152;
            BLU=8'd108;
        end
        4235:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4236:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4237:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4238:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4239:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4240:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4241:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4242:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4243:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4244:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4245:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4246:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4247:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4248:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4249:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4250:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4251:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4252:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4253:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4254:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4255:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4256:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4257:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4258:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4259:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4260:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4261:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4262:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4263:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4264:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4265:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4266:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4267:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4268:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4269:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4270:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4271:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4272:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4273:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4274:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4275:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4276:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4277:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4278:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4279:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4280:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4281:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4282:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4283:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4284:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4285:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4286:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4287:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4288:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4289:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4290:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4291:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4292:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4293:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4294:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4295:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4296:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4297:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4298:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4299:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4300:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4301:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4302:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4303:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4304:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4305:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4306:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4307:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4308:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4309:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4310:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4311:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4312:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4313:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4314:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4315:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4316:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4317:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4318:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4319:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4320:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4321:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4322:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4323:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4324:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4325:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4326:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4327:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4328:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4329:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4330:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4331:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4332:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4333:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4334:
        begin
            RED=8'd139;
            GRN=8'd139;
            BLU=8'd123;
        end
        4335:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        4336:
        begin
            RED=8'd232;
            GRN=8'd222;
            BLU=8'd25;
        end
        4337:
        begin
            RED=8'd208;
            GRN=8'd200;
            BLU=8'd50;
        end
        4338:
        begin
            RED=8'd127;
            GRN=8'd129;
            BLU=8'd136;
        end
        4339:
        begin
            RED=8'd74;
            GRN=8'd82;
            BLU=8'd193;
        end
        4340:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4341:
        begin
            RED=8'd62;
            GRN=8'd70;
            BLU=8'd199;
        end
        4342:
        begin
            RED=8'd32;
            GRN=8'd37;
            BLU=8'd104;
        end
        4343:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4352:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4353:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4354:
        begin
            RED=8'd21;
            GRN=8'd23;
            BLU=8'd68;
        end
        4355:
        begin
            RED=8'd57;
            GRN=8'd65;
            BLU=8'd184;
        end
        4356:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4357:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4358:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4359:
        begin
            RED=8'd78;
            GRN=8'd85;
            BLU=8'd188;
        end
        4360:
        begin
            RED=8'd132;
            GRN=8'd133;
            BLU=8'd131;
        end
        4361:
        begin
            RED=8'd132;
            GRN=8'd133;
            BLU=8'd131;
        end
        4362:
        begin
            RED=8'd122;
            GRN=8'd124;
            BLU=8'd141;
        end
        4363:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4364:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4365:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4366:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4367:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4368:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4369:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4370:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4371:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4372:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4373:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4374:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4375:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4376:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4377:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4378:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4379:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4380:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4381:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4382:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4383:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4384:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4385:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4386:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4387:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4388:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4389:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4390:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4391:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4392:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4393:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4394:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4395:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4396:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4397:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4398:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4399:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4400:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4401:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4402:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4403:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4404:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4405:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4406:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4407:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4408:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4409:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4410:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4411:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4412:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4413:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4414:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4415:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4416:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4417:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4418:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4419:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4420:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4421:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4422:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4423:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4424:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4425:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4426:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4427:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4428:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4429:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4430:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4431:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4432:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4433:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4434:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4435:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4436:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4437:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4438:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4439:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4440:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4441:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4442:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4443:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4444:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4445:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4446:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4447:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4448:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4449:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4450:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4451:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4452:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4453:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4454:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4455:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4456:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4457:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4458:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4459:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4460:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4461:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4462:
        begin
            RED=8'd90;
            GRN=8'd96;
            BLU=8'd175;
        end
        4463:
        begin
            RED=8'd132;
            GRN=8'd133;
            BLU=8'd131;
        end
        4464:
        begin
            RED=8'd78;
            GRN=8'd85;
            BLU=8'd188;
        end
        4465:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4466:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4467:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4468:
        begin
            RED=8'd59;
            GRN=8'd68;
            BLU=8'd191;
        end
        4469:
        begin
            RED=8'd30;
            GRN=8'd34;
            BLU=8'd95;
        end
        4470:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4471:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4480:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4481:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4482:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4483:
        begin
            RED=8'd6;
            GRN=8'd7;
            BLU=8'd19;
        end
        4484:
        begin
            RED=8'd30;
            GRN=8'd34;
            BLU=8'd96;
        end
        4485:
        begin
            RED=8'd57;
            GRN=8'd65;
            BLU=8'd183;
        end
        4486:
        begin
            RED=8'd62;
            GRN=8'd71;
            BLU=8'd200;
        end
        4487:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4488:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4489:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4490:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4491:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4492:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4493:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4494:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4495:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4496:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4497:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4498:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4499:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4500:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4501:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4502:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4503:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4504:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4505:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4506:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4507:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4508:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4509:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4510:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4511:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4512:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4513:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4514:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4515:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4516:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4517:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4518:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4519:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4520:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4521:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4522:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4523:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4524:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4525:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4526:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4527:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4528:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4529:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4530:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4531:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4532:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4533:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4534:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4535:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4536:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4537:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4538:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4539:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4540:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4541:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4542:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4543:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4544:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4545:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4546:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4547:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4548:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4549:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4550:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4551:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4552:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4553:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4554:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4555:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4556:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4557:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4558:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4559:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4560:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4561:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4562:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4563:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4564:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4565:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4566:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4567:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4568:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4569:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4570:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4571:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4572:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4573:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4574:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4575:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4576:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4577:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4578:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4579:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4580:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4581:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4582:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4583:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4584:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4585:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4586:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4587:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4588:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4589:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4590:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4591:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4592:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4593:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4594:
        begin
            RED=8'd57;
            GRN=8'd65;
            BLU=8'd185;
        end
        4595:
        begin
            RED=8'd30;
            GRN=8'd34;
            BLU=8'd96;
        end
        4596:
        begin
            RED=8'd12;
            GRN=8'd14;
            BLU=8'd40;
        end
        4597:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4598:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4599:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4608:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4609:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4610:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4611:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4612:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4613:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4614:
        begin
            RED=8'd21;
            GRN=8'd24;
            BLU=8'd69;
        end
        4615:
        begin
            RED=8'd33;
            GRN=8'd37;
            BLU=8'd106;
        end
        4616:
        begin
            RED=8'd58;
            GRN=8'd66;
            BLU=8'd188;
        end
        4617:
        begin
            RED=8'd58;
            GRN=8'd66;
            BLU=8'd188;
        end
        4618:
        begin
            RED=8'd62;
            GRN=8'd71;
            BLU=8'd201;
        end
        4619:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4620:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4621:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4622:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4623:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4624:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4625:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4626:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4627:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4628:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4629:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4630:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4631:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4632:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4633:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4634:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4635:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4636:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4637:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4638:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4639:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4640:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4641:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4642:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4643:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4644:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4645:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4646:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4647:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4648:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4649:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4650:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4651:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4652:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4653:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4654:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4655:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4656:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4657:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4658:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4659:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4660:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4661:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4662:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4663:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4664:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4665:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4666:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4667:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4668:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4669:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4670:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4671:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4672:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4673:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4674:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4675:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4676:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4677:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4678:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4679:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4680:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4681:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4682:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4683:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4684:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4685:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4686:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4687:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4688:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4689:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4690:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4691:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4692:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4693:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4694:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4695:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4696:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4697:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4698:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4699:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4700:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4701:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4702:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4703:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4704:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4705:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4706:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4707:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4708:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4709:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4710:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4711:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4712:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4713:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4714:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4715:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4716:
        begin
            RED=8'd63;
            GRN=8'd72;
            BLU=8'd204;
        end
        4717:
        begin
            RED=8'd62;
            GRN=8'd71;
            BLU=8'd201;
        end
        4718:
        begin
            RED=8'd58;
            GRN=8'd66;
            BLU=8'd188;
        end
        4719:
        begin
            RED=8'd58;
            GRN=8'd66;
            BLU=8'd188;
        end
        4720:
        begin
            RED=8'd33;
            GRN=8'd37;
            BLU=8'd106;
        end
        4721:
        begin
            RED=8'd26;
            GRN=8'd30;
            BLU=8'd84;
        end
        4722:
        begin
            RED=8'd2;
            GRN=8'd3;
            BLU=8'd8;
        end
        4723:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4724:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4725:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4726:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4727:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4736:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4737:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4738:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4739:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4740:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4741:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4742:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4743:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4744:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4745:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4746:
        begin
            RED=8'd40;
            GRN=8'd47;
            BLU=8'd132;
        end
        4747:
        begin
            RED=8'd56;
            GRN=8'd64;
            BLU=8'd183;
        end
        4748:
        begin
            RED=8'd27;
            GRN=8'd31;
            BLU=8'd89;
        end
        4749:
        begin
            RED=8'd46;
            GRN=8'd53;
            BLU=8'd149;
        end
        4750:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4751:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4752:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4753:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4754:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4755:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4756:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4757:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4758:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4759:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4760:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4761:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4762:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4763:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4764:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4765:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4766:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4767:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4768:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4769:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4770:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4771:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4772:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4773:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4774:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4775:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4776:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4777:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4778:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4779:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4780:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4781:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4782:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4783:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4784:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4785:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4786:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4787:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4788:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4789:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4790:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4791:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4792:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4793:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4794:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4795:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4796:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4797:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4798:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4799:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4800:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4801:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4802:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4803:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4804:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4805:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4806:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4807:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4808:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4809:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4810:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4811:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4812:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4813:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4814:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4815:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4816:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4817:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4818:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4819:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4820:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4821:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4822:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4823:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4824:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4825:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4826:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4827:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4828:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4829:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4830:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4831:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4832:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4833:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4834:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4835:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4836:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4837:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4838:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4839:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4840:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4841:
        begin
            RED=8'd60;
            GRN=8'd68;
            BLU=8'd194;
        end
        4842:
        begin
            RED=8'd46;
            GRN=8'd53;
            BLU=8'd149;
        end
        4843:
        begin
            RED=8'd27;
            GRN=8'd31;
            BLU=8'd89;
        end
        4844:
        begin
            RED=8'd27;
            GRN=8'd31;
            BLU=8'd89;
        end
        4845:
        begin
            RED=8'd22;
            GRN=8'd25;
            BLU=8'd71;
        end
        4846:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4847:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4848:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4849:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4850:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4851:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4852:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4853:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4854:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4855:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4864:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4865:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4866:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4867:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4868:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4869:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4870:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4871:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4872:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4873:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4874:
        begin
            RED=8'd23;
            GRN=8'd27;
            BLU=8'd77;
        end
        4875:
        begin
            RED=8'd41;
            GRN=8'd47;
            BLU=8'd134;
        end
        4876:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4877:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4878:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4879:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4880:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4881:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4882:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4883:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4884:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4885:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4886:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4887:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4888:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4889:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4890:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4891:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4892:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4893:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4894:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4895:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4896:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4897:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4898:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4899:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4900:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4901:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4902:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4903:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4904:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4905:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4906:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4907:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4908:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4909:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4910:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4911:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4912:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4913:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4914:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4916:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4917:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4918:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4919:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4920:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4921:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4922:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4923:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4924:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4925:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4926:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4927:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4928:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4929:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4930:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4931:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4932:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4933:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4934:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4935:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4936:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4937:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4938:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4939:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4940:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4941:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4942:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4943:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4944:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4945:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4946:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4947:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4948:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4949:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4950:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4951:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4952:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4953:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4954:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4955:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4956:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4957:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4958:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4959:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4960:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4961:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4962:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4963:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4964:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4965:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4966:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4967:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4968:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4969:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4970:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4971:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4972:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4973:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4974:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4975:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4976:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4977:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4978:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4980:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4981:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4982:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4983:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4992:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4993:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4994:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4995:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4996:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4997:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4998:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        4999:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5000:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5001:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5002:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5003:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5004:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5005:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5006:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5007:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5008:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5009:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5010:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5011:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5012:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5013:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5014:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5015:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5016:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5017:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5018:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5019:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5020:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5021:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5022:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5023:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5026:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5027:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5028:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5029:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5030:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5031:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5032:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5033:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5034:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5035:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5036:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5037:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5038:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5039:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5040:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5041:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5042:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5044:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5045:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5046:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5047:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5048:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5049:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5050:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5051:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5052:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5053:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5054:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5055:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5056:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5057:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5058:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5059:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5060:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5061:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5062:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5063:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5064:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5065:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5066:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5067:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5068:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5069:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5070:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5071:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5072:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5073:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5074:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5075:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5076:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5077:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5078:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5079:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5080:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5081:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5082:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5083:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5084:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5085:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5086:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5087:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5088:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5089:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5090:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5091:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5092:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5093:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5094:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5095:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5096:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5097:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5098:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5099:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5100:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5101:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5102:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5103:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5104:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5105:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5108:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5109:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5110:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        5111:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        default:
        begin
            RED=8'h00;
            GRN=8'h00;
            BLU=8'h00;
        end
     endcase
endmodule