`timescale 1ns / 1ps
module yellowBlock_40x40_rom(
    input  [5:0] x_idx,
    input  [5:0] y_idx,
    output reg [7:0] RED,
    output reg [7:0] GRN,
    output reg [7:0] BLU);
always @ (*)
    case ({y_idx,x_idx})
        0:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        3:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        4:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        5:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        6:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        7:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        8:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        9:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        10:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        11:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        12:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        13:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        14:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        15:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        16:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        17:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        18:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        19:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        20:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        21:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        22:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        23:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        24:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        25:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        26:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        27:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        28:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        29:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        30:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        31:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        32:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        33:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        34:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        35:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        36:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        37:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        38:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        39:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        64:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        65:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        66:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        67:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        68:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        69:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        70:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        71:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        72:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        73:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        74:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        75:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        76:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        77:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        78:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        79:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        80:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        81:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        82:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        83:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        84:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        85:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        86:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        87:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        88:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        89:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        90:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        91:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        92:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        93:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        94:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        95:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        96:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        97:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        98:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        99:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        100:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        101:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        102:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        103:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        128:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        129:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        130:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        131:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        132:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        133:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        134:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        135:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        136:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        137:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        138:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        139:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        140:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        141:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        142:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        143:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        144:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        145:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        146:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        147:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        148:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        149:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        150:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        151:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        152:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        153:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        154:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        155:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        156:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        157:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        158:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        159:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        160:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        161:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        162:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        163:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        164:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        165:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        166:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        167:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        192:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        193:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        194:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        195:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        196:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        197:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        198:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        199:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        200:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        201:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        202:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        203:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        204:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        205:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        206:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        207:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        208:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        209:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        210:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        211:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        212:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        213:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        214:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        215:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        216:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        217:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        218:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        219:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        220:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        221:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        222:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        223:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        224:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        225:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        226:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        227:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        228:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        229:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        230:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        231:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        256:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        257:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        258:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        259:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        260:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        261:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        262:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        263:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        264:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        265:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        266:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        267:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        268:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        269:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        270:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        271:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        272:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        273:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        274:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        275:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        276:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        277:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        278:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        279:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        280:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        281:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        282:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        283:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        284:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        285:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        286:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        287:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        288:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        289:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        290:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        291:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        292:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        293:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        294:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        295:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        320:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        321:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        322:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        323:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        324:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        325:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        326:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        327:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        328:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        329:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        330:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        331:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        332:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        333:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        334:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        335:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        336:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        337:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        338:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        339:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        340:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        341:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        342:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        343:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        344:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        345:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        346:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        347:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        348:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        349:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        350:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        351:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        352:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        353:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        354:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        355:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        356:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        357:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        358:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        359:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        384:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        385:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        386:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        387:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        388:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        389:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        390:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        391:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        392:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        393:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        394:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        395:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        396:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        397:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        398:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        399:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        400:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        401:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        402:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        403:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        404:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        405:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        406:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        407:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        408:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        409:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        410:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        411:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        412:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        413:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        414:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        415:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        416:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        417:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        418:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        419:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        420:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        421:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        422:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        423:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        448:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        449:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        450:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        451:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        452:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        453:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        454:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        455:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        456:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        457:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        458:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        459:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        460:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        461:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        462:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        463:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        464:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        465:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        466:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        467:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        468:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        469:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        470:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        471:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        472:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        473:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        474:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        475:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        476:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        477:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        478:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        479:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        480:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        481:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        482:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        483:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        484:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        485:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        486:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        487:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        512:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        513:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        514:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        515:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        516:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        517:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        518:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        519:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        520:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        521:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        522:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        523:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        524:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        525:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        526:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        527:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        528:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        529:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        530:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        531:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        532:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        533:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        534:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        535:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        536:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        537:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        538:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        539:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        540:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        541:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        542:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        543:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        544:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        545:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        546:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        547:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        548:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        549:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        550:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        551:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        576:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        577:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        578:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        579:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        580:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        581:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        582:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        583:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        584:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        585:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        586:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        587:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        588:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        589:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        590:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        591:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        592:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        593:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        594:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        595:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        596:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        597:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        598:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        599:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        600:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        601:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        602:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        603:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        604:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        605:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        606:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        607:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        608:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        609:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        610:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        611:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        612:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        613:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        614:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        615:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        640:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        641:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        642:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        643:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        644:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        645:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        646:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        647:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        648:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        649:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        650:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        651:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        652:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        653:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        654:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        655:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        656:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        657:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        658:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        659:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        660:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        661:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        662:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        663:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        664:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        665:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        666:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        667:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        668:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        669:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        670:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        671:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        672:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        673:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        674:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        675:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        676:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        677:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        678:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        679:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        704:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        705:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        706:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        707:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        708:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        709:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        710:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        711:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        712:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        713:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        714:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        715:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        716:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        717:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        718:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        719:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        720:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        721:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        722:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        723:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        724:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        725:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        726:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        727:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        728:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        729:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        730:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        731:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        732:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        733:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        734:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        735:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        736:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        737:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        738:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        739:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        740:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        741:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        742:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        743:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        768:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        769:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        770:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        771:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        772:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        773:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        774:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        775:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        776:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        777:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        778:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        779:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        780:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        781:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        782:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        783:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        784:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        785:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        786:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        787:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        788:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        789:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        790:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        791:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        792:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        793:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        794:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        795:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        796:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        797:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        798:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        799:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        800:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        801:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        802:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        803:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        804:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        805:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        806:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        807:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        832:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        833:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        834:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        835:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        836:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        837:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        838:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        839:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        840:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        841:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        842:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        843:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        844:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        845:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        846:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        847:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        848:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        849:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        850:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        851:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        852:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        853:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        854:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        855:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        856:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        857:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        858:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        859:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        860:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        861:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        862:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        863:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        864:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        865:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        866:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        867:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        868:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        869:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        870:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        871:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        896:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        897:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        898:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        899:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        900:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        901:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        902:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        903:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        904:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        905:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        906:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        907:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        908:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        909:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        910:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        911:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        912:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        913:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        914:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        915:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        916:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        917:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        918:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        919:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        920:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        921:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        922:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        923:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        924:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        925:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        926:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        927:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        928:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        929:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        930:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        931:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        932:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        933:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        934:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        935:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        960:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        961:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        962:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        963:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        964:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        965:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        966:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        967:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        968:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        969:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        970:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        971:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        972:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        973:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        974:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        975:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        976:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        977:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        978:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        979:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        980:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        981:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        982:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        983:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        984:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        985:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        986:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        987:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        988:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        989:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        990:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        991:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        992:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        993:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        994:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        995:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        996:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        997:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        998:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        999:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1024:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1025:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1026:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1027:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1028:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1029:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1030:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1031:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1032:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1033:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1034:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1035:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1036:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1037:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1038:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1039:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1040:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1041:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1042:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1043:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1044:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1045:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1046:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1047:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1048:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1049:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1050:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1051:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1052:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1053:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1054:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1055:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1056:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1057:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1058:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1059:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1060:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1061:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1062:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1063:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1088:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1089:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1090:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1091:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1092:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1093:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1094:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1095:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1096:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1097:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1098:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1099:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1100:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1101:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1102:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1103:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1104:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1105:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1106:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1107:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1108:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1109:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1110:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1111:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1112:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1113:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1114:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1115:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1116:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1117:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1118:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1119:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1120:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1121:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1122:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1123:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1124:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1125:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1126:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1127:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1152:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1153:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1154:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1155:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1156:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1157:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1158:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1159:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1160:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1161:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1162:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1163:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1164:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1165:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1166:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1167:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1168:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1169:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1170:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1171:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1172:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1173:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1174:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1175:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1176:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1177:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1178:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1179:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1180:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1181:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1182:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1183:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1184:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1185:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1186:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1187:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1188:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1189:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1190:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1191:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1216:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1217:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1218:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1219:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1220:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1221:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1222:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1223:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1224:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1225:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1226:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1227:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1228:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1229:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1230:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1231:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1232:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1233:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1234:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1235:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1236:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1237:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1238:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1239:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1240:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1241:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1242:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1243:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1244:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1245:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1246:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1247:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1248:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1249:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1250:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1251:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1252:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1253:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1254:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1255:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1280:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1281:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1282:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1283:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1284:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1285:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1286:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1287:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1288:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1289:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1290:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1291:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1292:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1293:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1294:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1295:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1296:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1297:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1298:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1299:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1300:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1301:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1302:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1303:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1304:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1305:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1306:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1307:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1308:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1309:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1310:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1311:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1312:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1313:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1314:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1315:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1316:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1317:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1318:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1319:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1344:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1345:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1346:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1347:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1348:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1349:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1350:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1351:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1352:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1353:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1354:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1355:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1356:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1357:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1358:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1359:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1360:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1361:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1362:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1363:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1364:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1365:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1366:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1367:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1368:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1369:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1370:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1371:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1372:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1373:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1374:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1375:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1376:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1377:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1378:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1379:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1380:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1381:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1382:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1383:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1408:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1409:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1410:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1411:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1412:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1413:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1414:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1415:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1416:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1417:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1418:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1419:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1420:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1421:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1422:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1423:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1424:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1425:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1426:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1427:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1428:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1429:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1430:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1431:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1432:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1433:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1434:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1435:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1436:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1437:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1438:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1439:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1440:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1441:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1442:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1443:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1444:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1445:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1446:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1447:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1472:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1473:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1474:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1475:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1476:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1477:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1478:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1479:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1480:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1481:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1482:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1483:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1484:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1485:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1486:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1487:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1488:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1489:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1490:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1491:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1492:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1493:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1494:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1495:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1496:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1497:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1498:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1499:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1500:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1501:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1502:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1503:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1504:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1505:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1506:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1507:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1508:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1509:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1510:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1511:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1536:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1537:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1538:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1539:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1540:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1541:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1542:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1543:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1544:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1545:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1546:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1547:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1548:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1549:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1550:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1551:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1552:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1553:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1554:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1555:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1556:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1557:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1558:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1559:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1560:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1561:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1562:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1563:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1564:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1565:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1566:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1567:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1568:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1569:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1570:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1571:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1572:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1573:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1574:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1575:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1600:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1601:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1602:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1603:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1604:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1605:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1606:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1607:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1608:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1609:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1610:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1611:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1612:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1613:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1614:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1615:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1616:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1617:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1618:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1619:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1620:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1621:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1622:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1623:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1624:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1625:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1626:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1627:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1628:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1629:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1630:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1631:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1632:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1633:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1634:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1635:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1636:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1637:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1638:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1639:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1664:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1665:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1666:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1667:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1668:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1669:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1670:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1671:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1672:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1673:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1674:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1675:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1676:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1677:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1678:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1679:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1680:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1681:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1682:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1683:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1684:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1685:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1686:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1687:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1688:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1689:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1690:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1691:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1692:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1693:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1694:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1695:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1696:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1697:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1698:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1699:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1700:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1701:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1702:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1703:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1728:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1729:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1730:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1731:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1732:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1733:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1734:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1735:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1736:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1737:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1738:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1739:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1740:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1741:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1742:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1743:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1744:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1745:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1746:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1747:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1748:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1749:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1750:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1751:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1752:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1753:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1754:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1755:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1756:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1757:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1758:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1759:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1760:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1761:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1762:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1763:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1764:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1765:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1766:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1767:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1792:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1793:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1794:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1795:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1796:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1797:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1798:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1799:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1800:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1801:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1802:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1803:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1804:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1805:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1806:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1807:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1808:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1809:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1810:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1811:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1812:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1813:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1814:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1815:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1816:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1817:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1818:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1819:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1820:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1821:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1822:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1823:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1824:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1825:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1826:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1827:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1828:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1829:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1830:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1831:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1856:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1857:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1858:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1859:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1860:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1861:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1862:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1863:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1864:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1865:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1866:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1867:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1868:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1869:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1870:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1871:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1872:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1873:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1874:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1875:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1876:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1877:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1878:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1879:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1880:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1881:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1882:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1883:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1884:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1885:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1886:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1887:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1888:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1889:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1890:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1891:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1892:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1893:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1894:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1895:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1920:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1921:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1922:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1923:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1924:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1925:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1926:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1927:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1928:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1929:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1930:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1931:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1932:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1933:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1934:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1935:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1936:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1937:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1938:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1939:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1940:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1941:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1942:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1943:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1944:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1945:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1946:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1947:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1948:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1949:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1950:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1951:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1952:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1953:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1954:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1955:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1956:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1957:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1958:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1959:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1984:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1985:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1986:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1987:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1988:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1989:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1990:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1991:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1992:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1993:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1994:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1995:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1996:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1997:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1998:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        1999:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2000:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2001:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2002:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2003:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2004:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2005:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2006:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2007:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2008:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2009:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2010:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2011:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2012:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2013:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2014:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2015:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2016:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2017:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2018:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2019:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2020:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2021:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2022:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2023:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2048:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2049:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2050:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2051:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2052:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2053:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2054:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2055:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2056:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2057:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2058:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2059:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2060:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2061:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2062:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2063:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2064:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2065:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2066:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2067:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2068:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2069:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2070:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2071:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2072:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2073:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2074:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2075:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2076:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2077:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2078:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2079:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2080:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2081:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2082:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2083:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2084:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2085:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2086:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2087:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2112:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2113:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2114:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2115:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2116:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2117:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2118:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2119:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2120:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2121:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2122:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2123:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2124:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2125:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2126:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2127:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2128:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2129:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2130:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2131:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2132:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2133:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2134:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2135:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2136:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2137:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2138:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2139:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2140:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2141:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2142:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2143:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2144:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2145:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2146:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2147:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2148:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2149:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2150:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2151:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2176:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2177:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2178:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2179:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2180:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2181:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2182:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2183:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2184:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2185:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2186:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2187:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2188:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2189:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2190:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2191:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2192:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2193:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2194:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2195:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2196:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2197:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2198:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2199:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2200:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2201:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2202:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2203:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2204:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2205:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2206:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2207:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2208:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2209:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2210:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2211:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2212:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2213:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2214:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2215:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2240:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2241:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2242:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2243:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2244:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2245:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2246:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2247:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2248:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2249:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2250:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2251:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2252:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2253:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2254:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2255:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2256:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2257:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2258:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2259:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2260:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2261:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2262:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2263:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2264:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2265:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2266:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2267:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2268:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2269:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2270:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2271:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2272:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2273:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2274:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2275:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2276:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2277:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2278:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2279:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2304:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2305:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2306:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2307:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2308:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2309:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2310:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2311:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2312:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2313:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2314:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2315:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2316:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2317:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2318:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2319:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2320:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2321:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2322:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2323:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2324:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2325:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2326:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2327:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2328:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2329:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2330:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2331:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2332:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2333:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2334:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2335:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2336:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2337:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2338:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2339:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2340:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2341:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2342:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2343:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2368:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2369:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2370:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2371:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2372:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2373:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2374:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2375:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2376:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2377:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2378:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2379:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2380:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2381:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2382:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2383:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2384:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2385:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2386:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2387:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2388:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2389:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2390:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2391:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2392:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2393:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2394:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2395:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2396:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2397:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2398:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2399:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2400:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2401:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2402:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2403:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2404:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2405:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2406:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2407:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2432:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2433:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2434:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2435:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2436:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2437:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2438:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2439:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2440:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2441:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2442:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2443:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2444:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2445:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2446:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2447:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2448:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2449:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2450:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2451:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2452:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2453:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2454:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2455:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2456:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2457:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2458:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2459:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2460:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2461:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2462:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2463:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2464:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2465:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2466:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2467:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2468:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2469:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2470:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2471:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2496:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2497:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2498:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2499:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2500:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2501:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2502:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2503:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2504:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2505:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2506:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2507:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2508:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2509:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2510:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2511:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2512:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2513:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2514:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2515:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2516:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2517:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2518:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2519:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2520:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2521:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2522:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2523:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2524:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2525:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2526:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2527:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2528:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2529:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2530:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2531:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2532:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2533:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2534:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        2535:
        begin
            RED=8'd255;
            GRN=8'd255;
            BLU=8'd0;
        end
        default:
        begin
            RED=8'h00;
            GRN=8'h00;
            BLU=8'h00;
        end
     endcase
endmodule