`timescale 1ns / 1ps
module ball_20x20_mask_rom(
    input  [5:0] x_idx,
    input  [5:0] y_idx,
    output reg [1:0] exist);
always @ (*)
    case ({y_idx,x_idx})
        0:
        begin
            exist=1'b0;
        end
        1:
        begin
            exist=1'b0;
        end
        2:
        begin
            exist=1'b0;
        end
        3:
        begin
            exist=1'b1;
        end
        4:
        begin
            exist=1'b1;
        end
        5:
        begin
            exist=1'b1;
        end
        6:
        begin
            exist=1'b1;
        end
        7:
        begin
            exist=1'b1;
        end
        8:
        begin
            exist=1'b1;
        end
        9:
        begin
            exist=1'b1;
        end
        10:
        begin
            exist=1'b1;
        end
        11:
        begin
            exist=1'b1;
        end
        12:
        begin
            exist=1'b1;
        end
        13:
        begin
            exist=1'b1;
        end
        14:
        begin
            exist=1'b1;
        end
        15:
        begin
            exist=1'b0;
        end
        16:
        begin
            exist=1'b0;
        end
        17:
        begin
            exist=1'b0;
        end
        18:
        begin
            exist=1'b0;
        end
        19:
        begin
            exist=1'b0;
        end
        64:
        begin
            exist=1'b0;
        end
        65:
        begin
            exist=1'b0;
        end
        66:
        begin
            exist=1'b0;
        end
        67:
        begin
            exist=1'b1;
        end
        68:
        begin
            exist=1'b1;
        end
        69:
        begin
            exist=1'b1;
        end
        70:
        begin
            exist=1'b1;
        end
        71:
        begin
            exist=1'b1;
        end
        72:
        begin
            exist=1'b1;
        end
        73:
        begin
            exist=1'b1;
        end
        74:
        begin
            exist=1'b1;
        end
        75:
        begin
            exist=1'b1;
        end
        76:
        begin
            exist=1'b1;
        end
        77:
        begin
            exist=1'b1;
        end
        78:
        begin
            exist=1'b1;
        end
        79:
        begin
            exist=1'b1;
        end
        80:
        begin
            exist=1'b0;
        end
        81:
        begin
            exist=1'b0;
        end
        82:
        begin
            exist=1'b0;
        end
        83:
        begin
            exist=1'b0;
        end
        128:
        begin
            exist=1'b0;
        end
        129:
        begin
            exist=1'b1;
        end
        130:
        begin
            exist=1'b1;
        end
        131:
        begin
            exist=1'b1;
        end
        132:
        begin
            exist=1'b1;
        end
        133:
        begin
            exist=1'b1;
        end
        134:
        begin
            exist=1'b1;
        end
        135:
        begin
            exist=1'b1;
        end
        136:
        begin
            exist=1'b1;
        end
        137:
        begin
            exist=1'b1;
        end
        138:
        begin
            exist=1'b0;
        end
        139:
        begin
            exist=1'b1;
        end
        140:
        begin
            exist=1'b1;
        end
        141:
        begin
            exist=1'b1;
        end
        142:
        begin
            exist=1'b1;
        end
        143:
        begin
            exist=1'b1;
        end
        144:
        begin
            exist=1'b1;
        end
        145:
        begin
            exist=1'b0;
        end
        146:
        begin
            exist=1'b1;
        end
        147:
        begin
            exist=1'b0;
        end
        192:
        begin
            exist=1'b0;
        end
        193:
        begin
            exist=1'b1;
        end
        194:
        begin
            exist=1'b1;
        end
        195:
        begin
            exist=1'b1;
        end
        196:
        begin
            exist=1'b1;
        end
        197:
        begin
            exist=1'b1;
        end
        198:
        begin
            exist=1'b1;
        end
        199:
        begin
            exist=1'b0;
        end
        200:
        begin
            exist=1'b1;
        end
        201:
        begin
            exist=1'b1;
        end
        202:
        begin
            exist=1'b1;
        end
        203:
        begin
            exist=1'b1;
        end
        204:
        begin
            exist=1'b0;
        end
        205:
        begin
            exist=1'b1;
        end
        206:
        begin
            exist=1'b1;
        end
        207:
        begin
            exist=1'b1;
        end
        208:
        begin
            exist=1'b1;
        end
        209:
        begin
            exist=1'b1;
        end
        210:
        begin
            exist=1'b0;
        end
        211:
        begin
            exist=1'b0;
        end
        256:
        begin
            exist=1'b1;
        end
        257:
        begin
            exist=1'b1;
        end
        258:
        begin
            exist=1'b1;
        end
        259:
        begin
            exist=1'b1;
        end
        260:
        begin
            exist=1'b1;
        end
        261:
        begin
            exist=1'b0;
        end
        262:
        begin
            exist=1'b0;
        end
        263:
        begin
            exist=1'b1;
        end
        264:
        begin
            exist=1'b1;
        end
        265:
        begin
            exist=1'b1;
        end
        266:
        begin
            exist=1'b1;
        end
        267:
        begin
            exist=1'b1;
        end
        268:
        begin
            exist=1'b1;
        end
        269:
        begin
            exist=1'b0;
        end
        270:
        begin
            exist=1'b1;
        end
        271:
        begin
            exist=1'b1;
        end
        272:
        begin
            exist=1'b1;
        end
        273:
        begin
            exist=1'b1;
        end
        274:
        begin
            exist=1'b0;
        end
        275:
        begin
            exist=1'b0;
        end
        320:
        begin
            exist=1'b1;
        end
        321:
        begin
            exist=1'b1;
        end
        322:
        begin
            exist=1'b1;
        end
        323:
        begin
            exist=1'b0;
        end
        324:
        begin
            exist=1'b1;
        end
        325:
        begin
            exist=1'b0;
        end
        326:
        begin
            exist=1'b0;
        end
        327:
        begin
            exist=1'b0;
        end
        328:
        begin
            exist=1'b0;
        end
        329:
        begin
            exist=1'b0;
        end
        330:
        begin
            exist=1'b0;
        end
        331:
        begin
            exist=1'b0;
        end
        332:
        begin
            exist=1'b0;
        end
        333:
        begin
            exist=1'b0;
        end
        334:
        begin
            exist=1'b1;
        end
        335:
        begin
            exist=1'b0;
        end
        336:
        begin
            exist=1'b1;
        end
        337:
        begin
            exist=1'b1;
        end
        338:
        begin
            exist=1'b1;
        end
        339:
        begin
            exist=1'b0;
        end
        384:
        begin
            exist=1'b1;
        end
        385:
        begin
            exist=1'b1;
        end
        386:
        begin
            exist=1'b1;
        end
        387:
        begin
            exist=1'b1;
        end
        388:
        begin
            exist=1'b0;
        end
        389:
        begin
            exist=1'b0;
        end
        390:
        begin
            exist=1'b0;
        end
        391:
        begin
            exist=1'b0;
        end
        392:
        begin
            exist=1'b0;
        end
        393:
        begin
            exist=1'b0;
        end
        394:
        begin
            exist=1'b0;
        end
        395:
        begin
            exist=1'b0;
        end
        396:
        begin
            exist=1'b0;
        end
        397:
        begin
            exist=1'b0;
        end
        398:
        begin
            exist=1'b1;
        end
        399:
        begin
            exist=1'b1;
        end
        400:
        begin
            exist=1'b1;
        end
        401:
        begin
            exist=1'b1;
        end
        402:
        begin
            exist=1'b1;
        end
        403:
        begin
            exist=1'b0;
        end
        448:
        begin
            exist=1'b1;
        end
        449:
        begin
            exist=1'b1;
        end
        450:
        begin
            exist=1'b1;
        end
        451:
        begin
            exist=1'b0;
        end
        452:
        begin
            exist=1'b1;
        end
        453:
        begin
            exist=1'b0;
        end
        454:
        begin
            exist=1'b0;
        end
        455:
        begin
            exist=1'b0;
        end
        456:
        begin
            exist=1'b0;
        end
        457:
        begin
            exist=1'b0;
        end
        458:
        begin
            exist=1'b0;
        end
        459:
        begin
            exist=1'b0;
        end
        460:
        begin
            exist=1'b0;
        end
        461:
        begin
            exist=1'b0;
        end
        462:
        begin
            exist=1'b1;
        end
        463:
        begin
            exist=1'b1;
        end
        464:
        begin
            exist=1'b0;
        end
        465:
        begin
            exist=1'b1;
        end
        466:
        begin
            exist=1'b1;
        end
        467:
        begin
            exist=1'b1;
        end
        512:
        begin
            exist=1'b1;
        end
        513:
        begin
            exist=1'b1;
        end
        514:
        begin
            exist=1'b1;
        end
        515:
        begin
            exist=1'b0;
        end
        516:
        begin
            exist=1'b1;
        end
        517:
        begin
            exist=1'b0;
        end
        518:
        begin
            exist=1'b0;
        end
        519:
        begin
            exist=1'b0;
        end
        520:
        begin
            exist=1'b0;
        end
        521:
        begin
            exist=1'b0;
        end
        522:
        begin
            exist=1'b0;
        end
        523:
        begin
            exist=1'b0;
        end
        524:
        begin
            exist=1'b0;
        end
        525:
        begin
            exist=1'b0;
        end
        526:
        begin
            exist=1'b1;
        end
        527:
        begin
            exist=1'b1;
        end
        528:
        begin
            exist=1'b1;
        end
        529:
        begin
            exist=1'b1;
        end
        530:
        begin
            exist=1'b1;
        end
        531:
        begin
            exist=1'b1;
        end
        576:
        begin
            exist=1'b1;
        end
        577:
        begin
            exist=1'b1;
        end
        578:
        begin
            exist=1'b1;
        end
        579:
        begin
            exist=1'b1;
        end
        580:
        begin
            exist=1'b1;
        end
        581:
        begin
            exist=1'b0;
        end
        582:
        begin
            exist=1'b0;
        end
        583:
        begin
            exist=1'b0;
        end
        584:
        begin
            exist=1'b0;
        end
        585:
        begin
            exist=1'b0;
        end
        586:
        begin
            exist=1'b0;
        end
        587:
        begin
            exist=1'b0;
        end
        588:
        begin
            exist=1'b0;
        end
        589:
        begin
            exist=1'b0;
        end
        590:
        begin
            exist=1'b0;
        end
        591:
        begin
            exist=1'b0;
        end
        592:
        begin
            exist=1'b0;
        end
        593:
        begin
            exist=1'b0;
        end
        594:
        begin
            exist=1'b1;
        end
        595:
        begin
            exist=1'b1;
        end
        640:
        begin
            exist=1'b1;
        end
        641:
        begin
            exist=1'b1;
        end
        642:
        begin
            exist=1'b0;
        end
        643:
        begin
            exist=1'b1;
        end
        644:
        begin
            exist=1'b0;
        end
        645:
        begin
            exist=1'b0;
        end
        646:
        begin
            exist=1'b0;
        end
        647:
        begin
            exist=1'b0;
        end
        648:
        begin
            exist=1'b0;
        end
        649:
        begin
            exist=1'b0;
        end
        650:
        begin
            exist=1'b0;
        end
        651:
        begin
            exist=1'b0;
        end
        652:
        begin
            exist=1'b0;
        end
        653:
        begin
            exist=1'b0;
        end
        654:
        begin
            exist=1'b0;
        end
        655:
        begin
            exist=1'b0;
        end
        656:
        begin
            exist=1'b0;
        end
        657:
        begin
            exist=1'b0;
        end
        658:
        begin
            exist=1'b1;
        end
        659:
        begin
            exist=1'b1;
        end
        704:
        begin
            exist=1'b1;
        end
        705:
        begin
            exist=1'b1;
        end
        706:
        begin
            exist=1'b1;
        end
        707:
        begin
            exist=1'b1;
        end
        708:
        begin
            exist=1'b0;
        end
        709:
        begin
            exist=1'b0;
        end
        710:
        begin
            exist=1'b0;
        end
        711:
        begin
            exist=1'b0;
        end
        712:
        begin
            exist=1'b0;
        end
        713:
        begin
            exist=1'b0;
        end
        714:
        begin
            exist=1'b0;
        end
        715:
        begin
            exist=1'b0;
        end
        716:
        begin
            exist=1'b0;
        end
        717:
        begin
            exist=1'b0;
        end
        718:
        begin
            exist=1'b0;
        end
        719:
        begin
            exist=1'b0;
        end
        720:
        begin
            exist=1'b0;
        end
        721:
        begin
            exist=1'b0;
        end
        722:
        begin
            exist=1'b1;
        end
        723:
        begin
            exist=1'b1;
        end
        768:
        begin
            exist=1'b1;
        end
        769:
        begin
            exist=1'b1;
        end
        770:
        begin
            exist=1'b1;
        end
        771:
        begin
            exist=1'b1;
        end
        772:
        begin
            exist=1'b0;
        end
        773:
        begin
            exist=1'b0;
        end
        774:
        begin
            exist=1'b0;
        end
        775:
        begin
            exist=1'b0;
        end
        776:
        begin
            exist=1'b0;
        end
        777:
        begin
            exist=1'b0;
        end
        778:
        begin
            exist=1'b0;
        end
        779:
        begin
            exist=1'b0;
        end
        780:
        begin
            exist=1'b0;
        end
        781:
        begin
            exist=1'b0;
        end
        782:
        begin
            exist=1'b0;
        end
        783:
        begin
            exist=1'b0;
        end
        784:
        begin
            exist=1'b0;
        end
        785:
        begin
            exist=1'b0;
        end
        786:
        begin
            exist=1'b1;
        end
        787:
        begin
            exist=1'b1;
        end
        832:
        begin
            exist=1'b1;
        end
        833:
        begin
            exist=1'b1;
        end
        834:
        begin
            exist=1'b1;
        end
        835:
        begin
            exist=1'b1;
        end
        836:
        begin
            exist=1'b1;
        end
        837:
        begin
            exist=1'b0;
        end
        838:
        begin
            exist=1'b0;
        end
        839:
        begin
            exist=1'b0;
        end
        840:
        begin
            exist=1'b0;
        end
        841:
        begin
            exist=1'b0;
        end
        842:
        begin
            exist=1'b0;
        end
        843:
        begin
            exist=1'b0;
        end
        844:
        begin
            exist=1'b0;
        end
        845:
        begin
            exist=1'b0;
        end
        846:
        begin
            exist=1'b0;
        end
        847:
        begin
            exist=1'b0;
        end
        848:
        begin
            exist=1'b0;
        end
        849:
        begin
            exist=1'b1;
        end
        850:
        begin
            exist=1'b1;
        end
        851:
        begin
            exist=1'b1;
        end
        896:
        begin
            exist=1'b1;
        end
        897:
        begin
            exist=1'b1;
        end
        898:
        begin
            exist=1'b1;
        end
        899:
        begin
            exist=1'b1;
        end
        900:
        begin
            exist=1'b0;
        end
        901:
        begin
            exist=1'b0;
        end
        902:
        begin
            exist=1'b0;
        end
        903:
        begin
            exist=1'b0;
        end
        904:
        begin
            exist=1'b0;
        end
        905:
        begin
            exist=1'b0;
        end
        906:
        begin
            exist=1'b0;
        end
        907:
        begin
            exist=1'b0;
        end
        908:
        begin
            exist=1'b0;
        end
        909:
        begin
            exist=1'b0;
        end
        910:
        begin
            exist=1'b1;
        end
        911:
        begin
            exist=1'b0;
        end
        912:
        begin
            exist=1'b1;
        end
        913:
        begin
            exist=1'b1;
        end
        914:
        begin
            exist=1'b1;
        end
        915:
        begin
            exist=1'b0;
        end
        960:
        begin
            exist=1'b1;
        end
        961:
        begin
            exist=1'b1;
        end
        962:
        begin
            exist=1'b1;
        end
        963:
        begin
            exist=1'b1;
        end
        964:
        begin
            exist=1'b1;
        end
        965:
        begin
            exist=1'b0;
        end
        966:
        begin
            exist=1'b0;
        end
        967:
        begin
            exist=1'b0;
        end
        968:
        begin
            exist=1'b0;
        end
        969:
        begin
            exist=1'b0;
        end
        970:
        begin
            exist=1'b0;
        end
        971:
        begin
            exist=1'b0;
        end
        972:
        begin
            exist=1'b0;
        end
        973:
        begin
            exist=1'b0;
        end
        974:
        begin
            exist=1'b0;
        end
        975:
        begin
            exist=1'b1;
        end
        976:
        begin
            exist=1'b1;
        end
        977:
        begin
            exist=1'b1;
        end
        978:
        begin
            exist=1'b0;
        end
        979:
        begin
            exist=1'b0;
        end
        1024:
        begin
            exist=1'b0;
        end
        1025:
        begin
            exist=1'b0;
        end
        1026:
        begin
            exist=1'b1;
        end
        1027:
        begin
            exist=1'b1;
        end
        1028:
        begin
            exist=1'b1;
        end
        1029:
        begin
            exist=1'b0;
        end
        1030:
        begin
            exist=1'b0;
        end
        1031:
        begin
            exist=1'b0;
        end
        1032:
        begin
            exist=1'b0;
        end
        1033:
        begin
            exist=1'b0;
        end
        1034:
        begin
            exist=1'b0;
        end
        1035:
        begin
            exist=1'b0;
        end
        1036:
        begin
            exist=1'b0;
        end
        1037:
        begin
            exist=1'b0;
        end
        1038:
        begin
            exist=1'b1;
        end
        1039:
        begin
            exist=1'b1;
        end
        1040:
        begin
            exist=1'b1;
        end
        1041:
        begin
            exist=1'b1;
        end
        1042:
        begin
            exist=1'b0;
        end
        1043:
        begin
            exist=1'b0;
        end
        1088:
        begin
            exist=1'b1;
        end
        1089:
        begin
            exist=1'b0;
        end
        1090:
        begin
            exist=1'b1;
        end
        1091:
        begin
            exist=1'b1;
        end
        1092:
        begin
            exist=1'b1;
        end
        1093:
        begin
            exist=1'b1;
        end
        1094:
        begin
            exist=1'b0;
        end
        1095:
        begin
            exist=1'b0;
        end
        1096:
        begin
            exist=1'b0;
        end
        1097:
        begin
            exist=1'b0;
        end
        1098:
        begin
            exist=1'b0;
        end
        1099:
        begin
            exist=1'b0;
        end
        1100:
        begin
            exist=1'b0;
        end
        1101:
        begin
            exist=1'b1;
        end
        1102:
        begin
            exist=1'b1;
        end
        1103:
        begin
            exist=1'b1;
        end
        1104:
        begin
            exist=1'b1;
        end
        1105:
        begin
            exist=1'b1;
        end
        1106:
        begin
            exist=1'b0;
        end
        1107:
        begin
            exist=1'b0;
        end
        1152:
        begin
            exist=1'b0;
        end
        1153:
        begin
            exist=1'b0;
        end
        1154:
        begin
            exist=1'b0;
        end
        1155:
        begin
            exist=1'b0;
        end
        1156:
        begin
            exist=1'b1;
        end
        1157:
        begin
            exist=1'b1;
        end
        1158:
        begin
            exist=1'b1;
        end
        1159:
        begin
            exist=1'b1;
        end
        1160:
        begin
            exist=1'b1;
        end
        1161:
        begin
            exist=1'b1;
        end
        1162:
        begin
            exist=1'b1;
        end
        1163:
        begin
            exist=1'b1;
        end
        1164:
        begin
            exist=1'b1;
        end
        1165:
        begin
            exist=1'b1;
        end
        1166:
        begin
            exist=1'b1;
        end
        1167:
        begin
            exist=1'b1;
        end
        1168:
        begin
            exist=1'b0;
        end
        1169:
        begin
            exist=1'b0;
        end
        1170:
        begin
            exist=1'b0;
        end
        1171:
        begin
            exist=1'b0;
        end
        1216:
        begin
            exist=1'b0;
        end
        1217:
        begin
            exist=1'b0;
        end
        1218:
        begin
            exist=1'b0;
        end
        1219:
        begin
            exist=1'b0;
        end
        1220:
        begin
            exist=1'b0;
        end
        1221:
        begin
            exist=1'b1;
        end
        1222:
        begin
            exist=1'b1;
        end
        1223:
        begin
            exist=1'b1;
        end
        1224:
        begin
            exist=1'b1;
        end
        1225:
        begin
            exist=1'b1;
        end
        1226:
        begin
            exist=1'b1;
        end
        1227:
        begin
            exist=1'b1;
        end
        1228:
        begin
            exist=1'b1;
        end
        1229:
        begin
            exist=1'b1;
        end
        1230:
        begin
            exist=1'b1;
        end
        1231:
        begin
            exist=1'b1;
        end
        1232:
        begin
            exist=1'b0;
        end
        1233:
        begin
            exist=1'b0;
        end
        1234:
        begin
            exist=1'b0;
        end
        1235:
        begin
            exist=1'b0;
        end
        default:
        begin
            exist=1'b0;
        end
     endcase
endmodule