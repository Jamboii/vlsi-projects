`timescale 1ns / 1ps
module ball_20x20_rom(
    input  [5:0] x_idx,
    input  [5:0] y_idx,
    output reg [7:0] RED,
    output reg [7:0] GRN,
    output reg [7:0] BLU);
always @ (*)
    case ({y_idx,x_idx})
        0:
        begin
            RED=8'd1;
            GRN=8'd0;
            BLU=8'd2;
        end
        1:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        2:
        begin
            RED=8'd1;
            GRN=8'd0;
            BLU=8'd5;
        end
        3:
        begin
            RED=8'd2;
            GRN=8'd1;
            BLU=8'd1;
        end
        4:
        begin
            RED=8'd1;
            GRN=8'd2;
            BLU=8'd2;
        end
        5:
        begin
            RED=8'd23;
            GRN=8'd22;
            BLU=8'd8;
        end
        6:
        begin
            RED=8'd107;
            GRN=8'd103;
            BLU=8'd21;
        end
        7:
        begin
            RED=8'd183;
            GRN=8'd173;
            BLU=8'd32;
        end
        8:
        begin
            RED=8'd244;
            GRN=8'd235;
            BLU=8'd7;
        end
        9:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd2;
        end
        10:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd5;
        end
        11:
        begin
            RED=8'd184;
            GRN=8'd175;
            BLU=8'd31;
        end
        12:
        begin
            RED=8'd123;
            GRN=8'd119;
            BLU=8'd23;
        end
        13:
        begin
            RED=8'd33;
            GRN=8'd29;
            BLU=8'd9;
        end
        14:
        begin
            RED=8'd3;
            GRN=8'd3;
            BLU=8'd1;
        end
        15:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd2;
        end
        16:
        begin
            RED=8'd1;
            GRN=8'd0;
            BLU=8'd2;
        end
        17:
        begin
            RED=8'd1;
            GRN=8'd1;
            BLU=8'd0;
        end
        18:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd3;
        end
        19:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        64:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        65:
        begin
            RED=8'd2;
            GRN=8'd0;
            BLU=8'd1;
        end
        66:
        begin
            RED=8'd3;
            GRN=8'd0;
            BLU=8'd1;
        end
        67:
        begin
            RED=8'd5;
            GRN=8'd4;
            BLU=8'd1;
        end
        68:
        begin
            RED=8'd129;
            GRN=8'd120;
            BLU=8'd27;
        end
        69:
        begin
            RED=8'd234;
            GRN=8'd225;
            BLU=8'd24;
        end
        70:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd6;
        end
        71:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd2;
        end
        72:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        73:
        begin
            RED=8'd252;
            GRN=8'd242;
            BLU=8'd3;
        end
        74:
        begin
            RED=8'd253;
            GRN=8'd243;
            BLU=8'd1;
        end
        75:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd3;
        end
        76:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd2;
        end
        77:
        begin
            RED=8'd241;
            GRN=8'd228;
            BLU=8'd18;
        end
        78:
        begin
            RED=8'd149;
            GRN=8'd142;
            BLU=8'd30;
        end
        79:
        begin
            RED=8'd14;
            GRN=8'd10;
            BLU=8'd3;
        end
        80:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd3;
        end
        81:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        82:
        begin
            RED=8'd2;
            GRN=8'd0;
            BLU=8'd0;
        end
        83:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        128:
        begin
            RED=8'd1;
            GRN=8'd0;
            BLU=8'd4;
        end
        129:
        begin
            RED=8'd3;
            GRN=8'd1;
            BLU=8'd1;
        end
        130:
        begin
            RED=8'd26;
            GRN=8'd26;
            BLU=8'd10;
        end
        131:
        begin
            RED=8'd168;
            GRN=8'd162;
            BLU=8'd29;
        end
        132:
        begin
            RED=8'd252;
            GRN=8'd242;
            BLU=8'd6;
        end
        133:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd2;
        end
        134:
        begin
            RED=8'd253;
            GRN=8'd243;
            BLU=8'd1;
        end
        135:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd3;
        end
        136:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd3;
        end
        137:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd2;
        end
        138:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        139:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd1;
        end
        140:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        141:
        begin
            RED=8'd253;
            GRN=8'd243;
            BLU=8'd2;
        end
        142:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd3;
        end
        143:
        begin
            RED=8'd208;
            GRN=8'd197;
            BLU=8'd26;
        end
        144:
        begin
            RED=8'd43;
            GRN=8'd41;
            BLU=8'd14;
        end
        145:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        146:
        begin
            RED=8'd1;
            GRN=8'd1;
            BLU=8'd2;
        end
        147:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        192:
        begin
            RED=8'd2;
            GRN=8'd1;
            BLU=8'd0;
        end
        193:
        begin
            RED=8'd8;
            GRN=8'd6;
            BLU=8'd2;
        end
        194:
        begin
            RED=8'd168;
            GRN=8'd162;
            BLU=8'd27;
        end
        195:
        begin
            RED=8'd254;
            GRN=8'd240;
            BLU=8'd7;
        end
        196:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd2;
        end
        197:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd3;
        end
        198:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd2;
        end
        199:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        200:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd1;
        end
        201:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        202:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd2;
        end
        203:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd2;
        end
        204:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        205:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        206:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd2;
        end
        207:
        begin
            RED=8'd254;
            GRN=8'd240;
            BLU=8'd4;
        end
        208:
        begin
            RED=8'd195;
            GRN=8'd184;
            BLU=8'd24;
        end
        209:
        begin
            RED=8'd19;
            GRN=8'd14;
            BLU=8'd5;
        end
        210:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd1;
        end
        211:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        256:
        begin
            RED=8'd1;
            GRN=8'd1;
            BLU=8'd1;
        end
        257:
        begin
            RED=8'd140;
            GRN=8'd131;
            BLU=8'd30;
        end
        258:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd3;
        end
        259:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd1;
        end
        260:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd3;
        end
        261:
        begin
            RED=8'd253;
            GRN=8'd243;
            BLU=8'd0;
        end
        262:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        263:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd1;
        end
        264:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        265:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        266:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd3;
        end
        267:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        268:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd1;
        end
        269:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        270:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        271:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd2;
        end
        272:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd4;
        end
        273:
        begin
            RED=8'd171;
            GRN=8'd162;
            BLU=8'd28;
        end
        274:
        begin
            RED=8'd2;
            GRN=8'd2;
            BLU=8'd0;
        end
        275:
        begin
            RED=8'd1;
            GRN=8'd0;
            BLU=8'd0;
        end
        320:
        begin
            RED=8'd32;
            GRN=8'd29;
            BLU=8'd9;
        end
        321:
        begin
            RED=8'd237;
            GRN=8'd227;
            BLU=8'd21;
        end
        322:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd2;
        end
        323:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        324:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd1;
        end
        325:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        326:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        327:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        328:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        329:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        330:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        331:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        332:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        333:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        334:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd1;
        end
        335:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        336:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd4;
        end
        337:
        begin
            RED=8'd248;
            GRN=8'd240;
            BLU=8'd18;
        end
        338:
        begin
            RED=8'd52;
            GRN=8'd48;
            BLU=8'd16;
        end
        339:
        begin
            RED=8'd1;
            GRN=8'd0;
            BLU=8'd1;
        end
        384:
        begin
            RED=8'd108;
            GRN=8'd103;
            BLU=8'd20;
        end
        385:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd3;
        end
        386:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd4;
        end
        387:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        388:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd0;
        end
        389:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        390:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        391:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        392:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        393:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        394:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        395:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        396:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        397:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        398:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        399:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd1;
        end
        400:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd1;
        end
        401:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd2;
        end
        402:
        begin
            RED=8'd141;
            GRN=8'd133;
            BLU=8'd21;
        end
        403:
        begin
            RED=8'd0;
            GRN=8'd2;
            BLU=8'd1;
        end
        448:
        begin
            RED=8'd175;
            GRN=8'd168;
            BLU=8'd34;
        end
        449:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd1;
        end
        450:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd1;
        end
        451:
        begin
            RED=8'd253;
            GRN=8'd243;
            BLU=8'd0;
        end
        452:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd4;
        end
        453:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        454:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        455:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        456:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        457:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        458:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        459:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        460:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        461:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        462:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd1;
        end
        463:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd3;
        end
        464:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        465:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd2;
        end
        466:
        begin
            RED=8'd210;
            GRN=8'd197;
            BLU=8'd31;
        end
        467:
        begin
            RED=8'd2;
            GRN=8'd4;
            BLU=8'd1;
        end
        512:
        begin
            RED=8'd221;
            GRN=8'd209;
            BLU=8'd18;
        end
        513:
        begin
            RED=8'd253;
            GRN=8'd243;
            BLU=8'd1;
        end
        514:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd3;
        end
        515:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd0;
        end
        516:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd2;
        end
        517:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        518:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        519:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        520:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        521:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        522:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        523:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        524:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        525:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        526:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        527:
        begin
            RED=8'd252;
            GRN=8'd242;
            BLU=8'd3;
        end
        528:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd1;
        end
        529:
        begin
            RED=8'd252;
            GRN=8'd243;
            BLU=8'd2;
        end
        530:
        begin
            RED=8'd245;
            GRN=8'd234;
            BLU=8'd17;
        end
        531:
        begin
            RED=8'd30;
            GRN=8'd28;
            BLU=8'd9;
        end
        576:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd4;
        end
        577:
        begin
            RED=8'd252;
            GRN=8'd243;
            BLU=8'd1;
        end
        578:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd1;
        end
        579:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd1;
        end
        580:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd1;
        end
        581:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        582:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        583:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        584:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        585:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        586:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        587:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        588:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        589:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        590:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        591:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        592:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        593:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        594:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd9;
        end
        595:
        begin
            RED=8'd35;
            GRN=8'd33;
            BLU=8'd7;
        end
        640:
        begin
            RED=8'd250;
            GRN=8'd240;
            BLU=8'd10;
        end
        641:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd2;
        end
        642:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd0;
        end
        643:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd1;
        end
        644:
        begin
            RED=8'd253;
            GRN=8'd243;
            BLU=8'd0;
        end
        645:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        646:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        647:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        648:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        649:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        650:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        651:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        652:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        653:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        654:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        655:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        656:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        657:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        658:
        begin
            RED=8'd252;
            GRN=8'd241;
            BLU=8'd10;
        end
        659:
        begin
            RED=8'd35;
            GRN=8'd33;
            BLU=8'd7;
        end
        704:
        begin
            RED=8'd181;
            GRN=8'd173;
            BLU=8'd27;
        end
        705:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd2;
        end
        706:
        begin
            RED=8'd255;
            GRN=8'd242;
            BLU=8'd1;
        end
        707:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        708:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        709:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        710:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        711:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        712:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        713:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        714:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        715:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        716:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        717:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        718:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        719:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        720:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        721:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        722:
        begin
            RED=8'd221;
            GRN=8'd213;
            BLU=8'd26;
        end
        723:
        begin
            RED=8'd14;
            GRN=8'd11;
            BLU=8'd3;
        end
        768:
        begin
            RED=8'd135;
            GRN=8'd130;
            BLU=8'd25;
        end
        769:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd1;
        end
        770:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd1;
        end
        771:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd2;
        end
        772:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd0;
        end
        773:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        774:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        775:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        776:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        777:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        778:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        779:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        780:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        781:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        782:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        783:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        784:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        785:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        786:
        begin
            RED=8'd168;
            GRN=8'd160;
            BLU=8'd23;
        end
        787:
        begin
            RED=8'd3;
            GRN=8'd2;
            BLU=8'd2;
        end
        832:
        begin
            RED=8'd72;
            GRN=8'd70;
            BLU=8'd16;
        end
        833:
        begin
            RED=8'd252;
            GRN=8'd241;
            BLU=8'd11;
        end
        834:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd1;
        end
        835:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd3;
        end
        836:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd1;
        end
        837:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        838:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        839:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        840:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        841:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        842:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        843:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        844:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        845:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        846:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd0;
        end
        847:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        848:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        849:
        begin
            RED=8'd252;
            GRN=8'd241;
            BLU=8'd6;
        end
        850:
        begin
            RED=8'd106;
            GRN=8'd100;
            BLU=8'd22;
        end
        851:
        begin
            RED=8'd1;
            GRN=8'd1;
            BLU=8'd1;
        end
        896:
        begin
            RED=8'd6;
            GRN=8'd5;
            BLU=8'd1;
        end
        897:
        begin
            RED=8'd189;
            GRN=8'd182;
            BLU=8'd25;
        end
        898:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd2;
        end
        899:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd1;
        end
        900:
        begin
            RED=8'd252;
            GRN=8'd243;
            BLU=8'd0;
        end
        901:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        902:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        903:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        904:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        905:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        906:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        907:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        908:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        909:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        910:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd1;
        end
        911:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        912:
        begin
            RED=8'd253;
            GRN=8'd243;
            BLU=8'd1;
        end
        913:
        begin
            RED=8'd219;
            GRN=8'd210;
            BLU=8'd25;
        end
        914:
        begin
            RED=8'd9;
            GRN=8'd7;
            BLU=8'd2;
        end
        915:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        960:
        begin
            RED=8'd1;
            GRN=8'd1;
            BLU=8'd1;
        end
        961:
        begin
            RED=8'd49;
            GRN=8'd48;
            BLU=8'd14;
        end
        962:
        begin
            RED=8'd231;
            GRN=8'd221;
            BLU=8'd21;
        end
        963:
        begin
            RED=8'd255;
            GRN=8'd241;
            BLU=8'd2;
        end
        964:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd1;
        end
        965:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        966:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        967:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        968:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        969:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        970:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        971:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        972:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        973:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        974:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        975:
        begin
            RED=8'd255;
            GRN=8'd240;
            BLU=8'd1;
        end
        976:
        begin
            RED=8'd242;
            GRN=8'd230;
            BLU=8'd17;
        end
        977:
        begin
            RED=8'd70;
            GRN=8'd72;
            BLU=8'd17;
        end
        978:
        begin
            RED=8'd1;
            GRN=8'd0;
            BLU=8'd1;
        end
        979:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1024:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd3;
        end
        1025:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd4;
        end
        1026:
        begin
            RED=8'd74;
            GRN=8'd72;
            BLU=8'd17;
        end
        1027:
        begin
            RED=8'd246;
            GRN=8'd236;
            BLU=8'd20;
        end
        1028:
        begin
            RED=8'd255;
            GRN=8'd240;
            BLU=8'd3;
        end
        1029:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1030:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1031:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1032:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1033:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1034:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1035:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1036:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1037:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1038:
        begin
            RED=8'd253;
            GRN=8'd242;
            BLU=8'd1;
        end
        1039:
        begin
            RED=8'd249;
            GRN=8'd239;
            BLU=8'd17;
        end
        1040:
        begin
            RED=8'd106;
            GRN=8'd99;
            BLU=8'd24;
        end
        1041:
        begin
            RED=8'd2;
            GRN=8'd1;
            BLU=8'd2;
        end
        1042:
        begin
            RED=8'd1;
            GRN=8'd0;
            BLU=8'd2;
        end
        1043:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1088:
        begin
            RED=8'd1;
            GRN=8'd2;
            BLU=8'd1;
        end
        1089:
        begin
            RED=8'd1;
            GRN=8'd0;
            BLU=8'd2;
        end
        1090:
        begin
            RED=8'd2;
            GRN=8'd1;
            BLU=8'd1;
        end
        1091:
        begin
            RED=8'd57;
            GRN=8'd55;
            BLU=8'd16;
        end
        1092:
        begin
            RED=8'd227;
            GRN=8'd214;
            BLU=8'd26;
        end
        1093:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd4;
        end
        1094:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1095:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1096:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1097:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1098:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1099:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1100:
        begin
            RED=8'd254;
            GRN=8'd242;
            BLU=8'd0;
        end
        1101:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd3;
        end
        1102:
        begin
            RED=8'd237;
            GRN=8'd226;
            BLU=8'd23;
        end
        1103:
        begin
            RED=8'd77;
            GRN=8'd73;
            BLU=8'd20;
        end
        1104:
        begin
            RED=8'd3;
            GRN=8'd2;
            BLU=8'd1;
        end
        1105:
        begin
            RED=8'd1;
            GRN=8'd1;
            BLU=8'd1;
        end
        1106:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1107:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1152:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1153:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1154:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1155:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1156:
        begin
            RED=8'd14;
            GRN=8'd11;
            BLU=8'd3;
        end
        1157:
        begin
            RED=8'd113;
            GRN=8'd110;
            BLU=8'd24;
        end
        1158:
        begin
            RED=8'd212;
            GRN=8'd205;
            BLU=8'd31;
        end
        1159:
        begin
            RED=8'd252;
            GRN=8'd240;
            BLU=8'd12;
        end
        1160:
        begin
            RED=8'd254;
            GRN=8'd241;
            BLU=8'd4;
        end
        1161:
        begin
            RED=8'd251;
            GRN=8'd243;
            BLU=8'd4;
        end
        1162:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd4;
        end
        1163:
        begin
            RED=8'd253;
            GRN=8'd241;
            BLU=8'd12;
        end
        1164:
        begin
            RED=8'd223;
            GRN=8'd215;
            BLU=8'd28;
        end
        1165:
        begin
            RED=8'd126;
            GRN=8'd121;
            BLU=8'd24;
        end
        1166:
        begin
            RED=8'd22;
            GRN=8'd23;
            BLU=8'd8;
        end
        1167:
        begin
            RED=8'd2;
            GRN=8'd1;
            BLU=8'd5;
        end
        1168:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd2;
        end
        1169:
        begin
            RED=8'd0;
            GRN=8'd1;
            BLU=8'd0;
        end
        1170:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        1171:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1216:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1217:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1218:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1219:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1220:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1221:
        begin
            RED=8'd2;
            GRN=8'd1;
            BLU=8'd2;
        end
        1222:
        begin
            RED=8'd7;
            GRN=8'd5;
            BLU=8'd1;
        end
        1223:
        begin
            RED=8'd41;
            GRN=8'd39;
            BLU=8'd10;
        end
        1224:
        begin
            RED=8'd102;
            GRN=8'd99;
            BLU=8'd26;
        end
        1225:
        begin
            RED=8'd114;
            GRN=8'd106;
            BLU=8'd29;
        end
        1226:
        begin
            RED=8'd110;
            GRN=8'd106;
            BLU=8'd29;
        end
        1227:
        begin
            RED=8'd44;
            GRN=8'd40;
            BLU=8'd10;
        end
        1228:
        begin
            RED=8'd11;
            GRN=8'd9;
            BLU=8'd3;
        end
        1229:
        begin
            RED=8'd2;
            GRN=8'd1;
            BLU=8'd2;
        end
        1230:
        begin
            RED=8'd2;
            GRN=8'd1;
            BLU=8'd4;
        end
        1231:
        begin
            RED=8'd1;
            GRN=8'd1;
            BLU=8'd3;
        end
        1232:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        1233:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        1234:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd1;
        end
        1235:
        begin
            RED=8'd0;
            GRN=8'd0;
            BLU=8'd0;
        end
        default:
        begin
            RED=8'h00;
            GRN=8'h00;
            BLU=8'h00;
        end
     endcase
endmodule